magic
tech sky130A
magscale 1 2
timestamp 1681267127
<< nwell >>
rect 201 1716 1145 1824
rect 133 1500 1193 1716
rect 133 1384 1019 1500
<< pwell >>
rect 207 1128 1089 1254
rect 33 992 1089 1128
rect 207 720 1089 992
rect 33 584 1089 720
rect 73 202 1089 584
<< mvnmos >>
rect 112 1018 212 1102
rect 112 610 212 694
rect 286 228 386 1228
rect 442 228 542 1228
rect 598 228 698 1228
rect 754 228 854 1228
rect 910 228 1010 1228
<< mvpmos >>
rect 252 1450 372 1650
rect 428 1450 548 1650
rect 604 1450 724 1650
rect 780 1450 900 1650
rect 974 1566 1074 1650
<< mvndiff >>
rect 233 1158 286 1228
rect 233 1124 241 1158
rect 275 1124 286 1158
rect 233 1102 286 1124
rect 59 1090 112 1102
rect 59 1056 67 1090
rect 101 1056 112 1090
rect 59 1018 112 1056
rect 212 1090 286 1102
rect 212 1056 241 1090
rect 275 1056 286 1090
rect 212 1022 286 1056
rect 212 1018 241 1022
rect 233 988 241 1018
rect 275 988 286 1022
rect 233 954 286 988
rect 233 920 241 954
rect 275 920 286 954
rect 233 886 286 920
rect 233 852 241 886
rect 275 852 286 886
rect 233 818 286 852
rect 233 784 241 818
rect 275 784 286 818
rect 233 750 286 784
rect 233 716 241 750
rect 275 716 286 750
rect 233 694 286 716
rect 59 682 112 694
rect 59 648 67 682
rect 101 648 112 682
rect 59 610 112 648
rect 212 682 286 694
rect 212 648 241 682
rect 275 648 286 682
rect 212 614 286 648
rect 212 610 241 614
rect 233 580 241 610
rect 275 580 286 614
rect 233 546 286 580
rect 233 512 241 546
rect 275 512 286 546
rect 233 478 286 512
rect 233 444 241 478
rect 275 444 286 478
rect 233 410 286 444
rect 233 376 241 410
rect 275 376 286 410
rect 233 342 286 376
rect 233 308 241 342
rect 275 308 286 342
rect 233 274 286 308
rect 233 240 241 274
rect 275 240 286 274
rect 233 228 286 240
rect 386 1158 442 1228
rect 386 1124 397 1158
rect 431 1124 442 1158
rect 386 1090 442 1124
rect 386 1056 397 1090
rect 431 1056 442 1090
rect 386 1022 442 1056
rect 386 988 397 1022
rect 431 988 442 1022
rect 386 954 442 988
rect 386 920 397 954
rect 431 920 442 954
rect 386 886 442 920
rect 386 852 397 886
rect 431 852 442 886
rect 386 818 442 852
rect 386 784 397 818
rect 431 784 442 818
rect 386 750 442 784
rect 386 716 397 750
rect 431 716 442 750
rect 386 682 442 716
rect 386 648 397 682
rect 431 648 442 682
rect 386 614 442 648
rect 386 580 397 614
rect 431 580 442 614
rect 386 546 442 580
rect 386 512 397 546
rect 431 512 442 546
rect 386 478 442 512
rect 386 444 397 478
rect 431 444 442 478
rect 386 410 442 444
rect 386 376 397 410
rect 431 376 442 410
rect 386 342 442 376
rect 386 308 397 342
rect 431 308 442 342
rect 386 274 442 308
rect 386 240 397 274
rect 431 240 442 274
rect 386 228 442 240
rect 542 1158 598 1228
rect 542 1124 553 1158
rect 587 1124 598 1158
rect 542 1090 598 1124
rect 542 1056 553 1090
rect 587 1056 598 1090
rect 542 1022 598 1056
rect 542 988 553 1022
rect 587 988 598 1022
rect 542 954 598 988
rect 542 920 553 954
rect 587 920 598 954
rect 542 886 598 920
rect 542 852 553 886
rect 587 852 598 886
rect 542 818 598 852
rect 542 784 553 818
rect 587 784 598 818
rect 542 750 598 784
rect 542 716 553 750
rect 587 716 598 750
rect 542 682 598 716
rect 542 648 553 682
rect 587 648 598 682
rect 542 614 598 648
rect 542 580 553 614
rect 587 580 598 614
rect 542 546 598 580
rect 542 512 553 546
rect 587 512 598 546
rect 542 478 598 512
rect 542 444 553 478
rect 587 444 598 478
rect 542 410 598 444
rect 542 376 553 410
rect 587 376 598 410
rect 542 342 598 376
rect 542 308 553 342
rect 587 308 598 342
rect 542 274 598 308
rect 542 240 553 274
rect 587 240 598 274
rect 542 228 598 240
rect 698 1158 754 1228
rect 698 1124 709 1158
rect 743 1124 754 1158
rect 698 1090 754 1124
rect 698 1056 709 1090
rect 743 1056 754 1090
rect 698 1022 754 1056
rect 698 988 709 1022
rect 743 988 754 1022
rect 698 954 754 988
rect 698 920 709 954
rect 743 920 754 954
rect 698 886 754 920
rect 698 852 709 886
rect 743 852 754 886
rect 698 818 754 852
rect 698 784 709 818
rect 743 784 754 818
rect 698 750 754 784
rect 698 716 709 750
rect 743 716 754 750
rect 698 682 754 716
rect 698 648 709 682
rect 743 648 754 682
rect 698 614 754 648
rect 698 580 709 614
rect 743 580 754 614
rect 698 546 754 580
rect 698 512 709 546
rect 743 512 754 546
rect 698 478 754 512
rect 698 444 709 478
rect 743 444 754 478
rect 698 410 754 444
rect 698 376 709 410
rect 743 376 754 410
rect 698 342 754 376
rect 698 308 709 342
rect 743 308 754 342
rect 698 274 754 308
rect 698 240 709 274
rect 743 240 754 274
rect 698 228 754 240
rect 854 1158 910 1228
rect 854 1124 865 1158
rect 899 1124 910 1158
rect 854 1090 910 1124
rect 854 1056 865 1090
rect 899 1056 910 1090
rect 854 1022 910 1056
rect 854 988 865 1022
rect 899 988 910 1022
rect 854 954 910 988
rect 854 920 865 954
rect 899 920 910 954
rect 854 886 910 920
rect 854 852 865 886
rect 899 852 910 886
rect 854 818 910 852
rect 854 784 865 818
rect 899 784 910 818
rect 854 750 910 784
rect 854 716 865 750
rect 899 716 910 750
rect 854 682 910 716
rect 854 648 865 682
rect 899 648 910 682
rect 854 614 910 648
rect 854 580 865 614
rect 899 580 910 614
rect 854 546 910 580
rect 854 512 865 546
rect 899 512 910 546
rect 854 478 910 512
rect 854 444 865 478
rect 899 444 910 478
rect 854 410 910 444
rect 854 376 865 410
rect 899 376 910 410
rect 854 342 910 376
rect 854 308 865 342
rect 899 308 910 342
rect 854 274 910 308
rect 854 240 865 274
rect 899 240 910 274
rect 854 228 910 240
rect 1010 1158 1063 1228
rect 1010 1124 1021 1158
rect 1055 1124 1063 1158
rect 1010 1090 1063 1124
rect 1010 1056 1021 1090
rect 1055 1056 1063 1090
rect 1010 1022 1063 1056
rect 1010 988 1021 1022
rect 1055 988 1063 1022
rect 1010 954 1063 988
rect 1010 920 1021 954
rect 1055 920 1063 954
rect 1010 886 1063 920
rect 1010 852 1021 886
rect 1055 852 1063 886
rect 1010 818 1063 852
rect 1010 784 1021 818
rect 1055 784 1063 818
rect 1010 750 1063 784
rect 1010 716 1021 750
rect 1055 716 1063 750
rect 1010 682 1063 716
rect 1010 648 1021 682
rect 1055 648 1063 682
rect 1010 614 1063 648
rect 1010 580 1021 614
rect 1055 580 1063 614
rect 1010 546 1063 580
rect 1010 512 1021 546
rect 1055 512 1063 546
rect 1010 478 1063 512
rect 1010 444 1021 478
rect 1055 444 1063 478
rect 1010 410 1063 444
rect 1010 376 1021 410
rect 1055 376 1063 410
rect 1010 342 1063 376
rect 1010 308 1021 342
rect 1055 308 1063 342
rect 1010 274 1063 308
rect 1010 240 1021 274
rect 1055 240 1063 274
rect 1010 228 1063 240
<< mvpdiff >>
rect 199 1638 252 1650
rect 199 1604 207 1638
rect 241 1604 252 1638
rect 199 1570 252 1604
rect 199 1536 207 1570
rect 241 1536 252 1570
rect 199 1502 252 1536
rect 199 1468 207 1502
rect 241 1468 252 1502
rect 199 1450 252 1468
rect 372 1638 428 1650
rect 372 1604 383 1638
rect 417 1604 428 1638
rect 372 1570 428 1604
rect 372 1536 383 1570
rect 417 1536 428 1570
rect 372 1502 428 1536
rect 372 1468 383 1502
rect 417 1468 428 1502
rect 372 1450 428 1468
rect 548 1638 604 1650
rect 548 1604 559 1638
rect 593 1604 604 1638
rect 548 1570 604 1604
rect 548 1536 559 1570
rect 593 1536 604 1570
rect 548 1502 604 1536
rect 548 1468 559 1502
rect 593 1468 604 1502
rect 548 1450 604 1468
rect 724 1638 780 1650
rect 724 1604 735 1638
rect 769 1604 780 1638
rect 724 1570 780 1604
rect 724 1536 735 1570
rect 769 1536 780 1570
rect 724 1502 780 1536
rect 724 1468 735 1502
rect 769 1468 780 1502
rect 724 1450 780 1468
rect 900 1638 974 1650
rect 900 1604 911 1638
rect 945 1604 974 1638
rect 900 1570 974 1604
rect 900 1536 911 1570
rect 945 1566 974 1570
rect 1074 1638 1127 1650
rect 1074 1604 1085 1638
rect 1119 1604 1127 1638
rect 1074 1566 1127 1604
rect 945 1536 953 1566
rect 900 1502 953 1536
rect 900 1468 911 1502
rect 945 1468 953 1502
rect 900 1450 953 1468
<< mvndiffc >>
rect 241 1124 275 1158
rect 67 1056 101 1090
rect 241 1056 275 1090
rect 241 988 275 1022
rect 241 920 275 954
rect 241 852 275 886
rect 241 784 275 818
rect 241 716 275 750
rect 67 648 101 682
rect 241 648 275 682
rect 241 580 275 614
rect 241 512 275 546
rect 241 444 275 478
rect 241 376 275 410
rect 241 308 275 342
rect 241 240 275 274
rect 397 1124 431 1158
rect 397 1056 431 1090
rect 397 988 431 1022
rect 397 920 431 954
rect 397 852 431 886
rect 397 784 431 818
rect 397 716 431 750
rect 397 648 431 682
rect 397 580 431 614
rect 397 512 431 546
rect 397 444 431 478
rect 397 376 431 410
rect 397 308 431 342
rect 397 240 431 274
rect 553 1124 587 1158
rect 553 1056 587 1090
rect 553 988 587 1022
rect 553 920 587 954
rect 553 852 587 886
rect 553 784 587 818
rect 553 716 587 750
rect 553 648 587 682
rect 553 580 587 614
rect 553 512 587 546
rect 553 444 587 478
rect 553 376 587 410
rect 553 308 587 342
rect 553 240 587 274
rect 709 1124 743 1158
rect 709 1056 743 1090
rect 709 988 743 1022
rect 709 920 743 954
rect 709 852 743 886
rect 709 784 743 818
rect 709 716 743 750
rect 709 648 743 682
rect 709 580 743 614
rect 709 512 743 546
rect 709 444 743 478
rect 709 376 743 410
rect 709 308 743 342
rect 709 240 743 274
rect 865 1124 899 1158
rect 865 1056 899 1090
rect 865 988 899 1022
rect 865 920 899 954
rect 865 852 899 886
rect 865 784 899 818
rect 865 716 899 750
rect 865 648 899 682
rect 865 580 899 614
rect 865 512 899 546
rect 865 444 899 478
rect 865 376 899 410
rect 865 308 899 342
rect 865 240 899 274
rect 1021 1124 1055 1158
rect 1021 1056 1055 1090
rect 1021 988 1055 1022
rect 1021 920 1055 954
rect 1021 852 1055 886
rect 1021 784 1055 818
rect 1021 716 1055 750
rect 1021 648 1055 682
rect 1021 580 1055 614
rect 1021 512 1055 546
rect 1021 444 1055 478
rect 1021 376 1055 410
rect 1021 308 1055 342
rect 1021 240 1055 274
<< mvpdiffc >>
rect 207 1604 241 1638
rect 207 1536 241 1570
rect 207 1468 241 1502
rect 383 1604 417 1638
rect 383 1536 417 1570
rect 383 1468 417 1502
rect 559 1604 593 1638
rect 559 1536 593 1570
rect 559 1468 593 1502
rect 735 1604 769 1638
rect 735 1536 769 1570
rect 735 1468 769 1502
rect 911 1604 945 1638
rect 911 1536 945 1570
rect 1085 1604 1119 1638
rect 911 1468 945 1502
<< psubdiff >>
rect 99 486 159 510
rect 99 452 112 486
rect 146 452 159 486
rect 99 386 159 452
rect 99 352 112 386
rect 146 352 159 386
rect 99 286 159 352
rect 99 252 112 286
rect 146 252 159 286
rect 99 228 159 252
<< mvnsubdiff >>
rect 267 1724 291 1758
rect 325 1724 364 1758
rect 398 1724 437 1758
rect 471 1724 510 1758
rect 544 1724 583 1758
rect 617 1724 656 1758
rect 690 1724 729 1758
rect 763 1724 802 1758
rect 836 1724 875 1758
rect 909 1724 948 1758
rect 982 1724 1021 1758
rect 1055 1724 1079 1758
<< psubdiffcont >>
rect 112 452 146 486
rect 112 352 146 386
rect 112 252 146 286
<< mvnsubdiffcont >>
rect 291 1724 325 1758
rect 364 1724 398 1758
rect 437 1724 471 1758
rect 510 1724 544 1758
rect 583 1724 617 1758
rect 656 1724 690 1758
rect 729 1724 763 1758
rect 802 1724 836 1758
rect 875 1724 909 1758
rect 948 1724 982 1758
rect 1021 1724 1055 1758
<< poly >>
rect 974 1517 1074 1566
rect 974 1483 1016 1517
rect 1050 1483 1074 1517
rect 252 1418 372 1450
rect 428 1418 548 1450
rect 252 1402 548 1418
rect 252 1368 268 1402
rect 302 1368 345 1402
rect 379 1368 422 1402
rect 456 1368 498 1402
rect 532 1368 548 1402
rect 252 1352 548 1368
rect 604 1418 724 1450
rect 780 1418 900 1450
rect 604 1402 900 1418
rect 604 1368 620 1402
rect 654 1368 696 1402
rect 730 1368 773 1402
rect 807 1368 850 1402
rect 884 1368 900 1402
rect 974 1449 1074 1483
rect 974 1415 1016 1449
rect 1050 1415 1074 1449
rect 974 1399 1074 1415
rect 604 1352 900 1368
rect 112 1271 212 1288
rect 112 1237 145 1271
rect 179 1237 212 1271
rect 112 1203 212 1237
rect 112 1169 145 1203
rect 179 1169 212 1203
rect 112 1102 212 1169
rect 112 863 212 880
rect 112 829 145 863
rect 179 829 212 863
rect 112 795 212 829
rect 112 761 145 795
rect 179 761 212 795
rect 112 694 212 761
rect 286 158 386 228
rect 286 124 319 158
rect 353 124 386 158
rect 286 90 386 124
rect 286 56 319 90
rect 353 56 386 90
rect 286 40 386 56
rect 442 158 542 228
rect 442 124 479 158
rect 513 124 542 158
rect 442 90 542 124
rect 442 56 479 90
rect 513 56 542 90
rect 442 40 542 56
rect 598 158 698 228
rect 598 124 635 158
rect 669 124 698 158
rect 598 90 698 124
rect 598 56 635 90
rect 669 56 698 90
rect 598 40 698 56
rect 754 158 854 228
rect 754 124 785 158
rect 819 124 854 158
rect 754 90 854 124
rect 754 56 785 90
rect 819 56 854 90
rect 754 40 854 56
rect 910 156 1010 228
rect 910 122 940 156
rect 974 122 1010 156
rect 910 88 1010 122
rect 910 54 940 88
rect 974 54 1010 88
rect 910 38 1010 54
<< polycont >>
rect 1016 1483 1050 1517
rect 268 1368 302 1402
rect 345 1368 379 1402
rect 422 1368 456 1402
rect 498 1368 532 1402
rect 620 1368 654 1402
rect 696 1368 730 1402
rect 773 1368 807 1402
rect 850 1368 884 1402
rect 1016 1415 1050 1449
rect 145 1237 179 1271
rect 145 1169 179 1203
rect 145 829 179 863
rect 145 761 179 795
rect 319 124 353 158
rect 319 56 353 90
rect 479 124 513 158
rect 479 56 513 90
rect 635 124 669 158
rect 635 56 669 90
rect 785 124 819 158
rect 785 56 819 90
rect 940 122 974 156
rect 940 54 974 88
<< locali >>
rect 267 1724 291 1758
rect 325 1724 326 1758
rect 360 1724 364 1758
rect 398 1724 402 1758
rect 436 1724 437 1758
rect 471 1724 478 1758
rect 544 1724 554 1758
rect 617 1724 630 1758
rect 690 1724 706 1758
rect 763 1724 782 1758
rect 836 1724 858 1758
rect 909 1724 934 1758
rect 982 1724 1011 1758
rect 1055 1724 1079 1758
rect 911 1679 945 1724
rect 207 1582 241 1604
rect 207 1510 241 1536
rect 207 1452 241 1468
rect 383 1582 417 1604
rect 383 1510 417 1536
rect 383 1452 417 1468
rect 559 1582 593 1604
rect 559 1510 593 1536
rect 559 1452 593 1468
rect 735 1582 769 1604
rect 735 1510 769 1536
rect 735 1452 769 1468
rect 911 1638 945 1645
rect 1047 1620 1085 1654
rect 911 1597 945 1604
rect 1085 1588 1119 1604
rect 911 1502 945 1536
rect 911 1452 945 1468
rect 996 1522 1011 1549
rect 1045 1522 1119 1549
rect 996 1517 1119 1522
rect 996 1484 1016 1517
rect 996 1450 1011 1484
rect 1050 1483 1119 1517
rect 1045 1450 1119 1483
rect 996 1449 1119 1450
rect 996 1415 1016 1449
rect 1050 1415 1119 1449
rect 252 1368 268 1402
rect 302 1368 345 1402
rect 379 1368 422 1402
rect 456 1368 498 1402
rect 532 1368 548 1402
rect 604 1368 620 1402
rect 654 1368 696 1402
rect 730 1368 773 1402
rect 807 1368 850 1402
rect 884 1400 900 1402
rect 884 1368 902 1400
rect 996 1399 1119 1415
rect 119 1299 154 1333
rect 188 1299 226 1333
rect 119 1271 225 1299
rect 119 1237 145 1271
rect 179 1237 225 1271
rect 119 1205 225 1237
rect 119 1203 203 1205
rect 119 1169 145 1203
rect 179 1169 203 1203
rect 309 1181 363 1368
rect 604 1356 902 1368
rect 604 1322 658 1356
rect 692 1322 748 1356
rect 782 1322 838 1356
rect 872 1322 902 1356
rect 604 1316 902 1322
rect 119 1153 203 1169
rect 241 1158 275 1174
rect 67 1090 158 1106
rect 101 1072 158 1090
rect 101 1056 192 1072
rect 67 1040 192 1056
rect 119 1034 192 1040
rect 119 1000 158 1034
rect 119 863 192 1000
rect 119 829 145 863
rect 179 829 192 863
rect 119 795 192 829
rect 119 761 145 795
rect 179 761 192 795
rect 119 745 192 761
rect 241 1092 275 1124
rect 309 1147 320 1181
rect 354 1147 363 1181
rect 309 1109 363 1147
rect 309 1075 320 1109
rect 354 1075 363 1109
rect 309 1074 363 1075
rect 397 1158 431 1174
rect 397 1090 431 1124
rect 241 1022 275 1056
rect 241 954 275 984
rect 241 886 275 910
rect 241 818 275 836
rect 241 750 275 761
rect 67 682 158 698
rect 101 664 158 682
rect 101 648 192 664
rect 67 632 192 648
rect 158 626 192 632
rect 241 682 275 686
rect 241 645 275 648
rect 241 570 275 580
rect 99 492 159 510
rect 241 495 275 512
rect 99 486 118 492
rect 99 452 112 486
rect 152 458 165 492
rect 146 452 165 458
rect 99 414 165 452
rect 99 386 118 414
rect 99 352 112 386
rect 152 380 165 414
rect 146 352 165 380
rect 99 336 165 352
rect 99 302 118 336
rect 152 302 165 336
rect 99 286 165 302
rect 99 252 112 286
rect 146 258 165 286
rect 99 228 118 252
rect 105 224 118 228
rect 152 224 165 258
rect 241 420 275 444
rect 241 345 275 376
rect 397 1022 431 1056
rect 397 954 431 972
rect 397 886 431 899
rect 397 818 431 826
rect 397 750 431 753
rect 397 714 431 716
rect 397 640 431 648
rect 397 566 431 580
rect 397 492 431 512
rect 397 418 431 444
rect 397 344 431 376
rect 241 274 275 308
rect 241 224 275 236
rect 311 309 320 343
rect 354 309 361 343
rect 311 271 361 309
rect 311 237 320 271
rect 354 237 361 271
rect 311 158 361 237
rect 397 274 431 308
rect 397 224 431 236
rect 553 1158 587 1174
rect 553 1090 587 1124
rect 553 1022 587 1056
rect 553 954 587 972
rect 553 886 587 899
rect 553 818 587 826
rect 553 750 587 753
rect 553 714 587 716
rect 553 640 587 648
rect 553 566 587 580
rect 553 492 587 512
rect 553 418 587 444
rect 553 344 587 376
rect 553 274 587 308
rect 553 224 587 236
rect 709 1158 743 1174
rect 709 1090 743 1124
rect 709 1022 743 1056
rect 709 954 743 972
rect 709 886 743 899
rect 709 818 743 826
rect 709 750 743 753
rect 709 714 743 716
rect 709 640 743 648
rect 709 566 743 580
rect 709 492 743 512
rect 709 418 743 444
rect 709 344 743 376
rect 709 274 743 308
rect 709 224 743 236
rect 865 1158 899 1174
rect 865 1090 899 1124
rect 865 1022 899 1056
rect 865 954 899 972
rect 865 886 899 899
rect 865 818 899 826
rect 865 750 899 753
rect 865 714 899 716
rect 865 640 899 648
rect 865 566 899 580
rect 865 492 899 512
rect 865 418 899 444
rect 865 344 899 376
rect 865 274 899 308
rect 865 224 899 236
rect 1021 1100 1055 1124
rect 1021 1026 1055 1056
rect 1021 954 1055 988
rect 1021 886 1055 918
rect 1021 818 1055 844
rect 1021 750 1055 770
rect 1021 682 1055 696
rect 1021 614 1055 622
rect 1021 546 1055 547
rect 1021 506 1055 512
rect 1021 410 1055 444
rect 1021 342 1055 376
rect 1021 274 1055 308
rect 1021 224 1055 240
rect 311 124 319 158
rect 353 124 361 158
rect 479 158 513 174
rect 311 90 361 124
rect 478 124 479 137
rect 635 158 669 174
rect 478 109 513 124
rect 634 124 635 137
rect 634 109 669 124
rect 311 56 319 90
rect 353 56 361 90
rect 311 40 361 56
rect 479 90 513 109
rect 479 40 513 56
rect 635 90 669 109
rect 635 40 669 56
rect 785 158 819 174
rect 785 90 819 124
rect 785 40 819 56
rect 940 156 974 172
rect 940 88 974 122
rect 940 38 974 54
<< viali >>
rect 326 1724 360 1758
rect 402 1724 436 1758
rect 478 1724 510 1758
rect 510 1724 512 1758
rect 554 1724 583 1758
rect 583 1724 588 1758
rect 630 1724 656 1758
rect 656 1724 664 1758
rect 706 1724 729 1758
rect 729 1724 740 1758
rect 782 1724 802 1758
rect 802 1724 816 1758
rect 858 1724 875 1758
rect 875 1724 892 1758
rect 934 1724 948 1758
rect 948 1724 968 1758
rect 1011 1724 1021 1758
rect 1021 1724 1045 1758
rect 207 1638 241 1654
rect 207 1620 241 1638
rect 207 1570 241 1582
rect 207 1548 241 1570
rect 207 1502 241 1510
rect 207 1476 241 1502
rect 383 1638 417 1654
rect 383 1620 417 1638
rect 383 1570 417 1582
rect 383 1548 417 1570
rect 383 1502 417 1510
rect 383 1476 417 1502
rect 559 1638 593 1654
rect 559 1620 593 1638
rect 559 1570 593 1582
rect 559 1548 593 1570
rect 559 1502 593 1510
rect 559 1476 593 1502
rect 735 1638 769 1654
rect 735 1620 769 1638
rect 735 1570 769 1582
rect 735 1548 769 1570
rect 735 1502 769 1510
rect 735 1476 769 1502
rect 911 1645 945 1679
rect 1013 1620 1047 1654
rect 1085 1638 1119 1654
rect 1085 1620 1119 1638
rect 911 1570 945 1597
rect 911 1563 945 1570
rect 1011 1522 1045 1556
rect 1011 1483 1016 1484
rect 1016 1483 1045 1484
rect 1011 1450 1045 1483
rect 154 1299 188 1333
rect 226 1299 260 1333
rect 658 1322 692 1356
rect 748 1322 782 1356
rect 838 1322 872 1356
rect 158 1072 192 1106
rect 158 1000 192 1034
rect 241 1090 275 1092
rect 241 1058 275 1090
rect 320 1147 354 1181
rect 320 1075 354 1109
rect 241 988 275 1018
rect 241 984 275 988
rect 241 920 275 944
rect 241 910 275 920
rect 241 852 275 870
rect 241 836 275 852
rect 241 784 275 795
rect 241 761 275 784
rect 241 716 275 720
rect 158 664 192 698
rect 158 592 192 626
rect 241 686 275 716
rect 241 614 275 645
rect 241 611 275 614
rect 241 546 275 570
rect 241 536 275 546
rect 118 486 152 492
rect 118 458 146 486
rect 146 458 152 486
rect 118 386 152 414
rect 118 380 146 386
rect 146 380 152 386
rect 118 302 152 336
rect 118 252 146 258
rect 146 252 152 258
rect 118 224 152 252
rect 241 478 275 495
rect 241 461 275 478
rect 241 410 275 420
rect 241 386 275 410
rect 241 342 275 345
rect 397 988 431 1006
rect 397 972 431 988
rect 397 920 431 933
rect 397 899 431 920
rect 397 852 431 860
rect 397 826 431 852
rect 397 784 431 787
rect 397 753 431 784
rect 397 682 431 714
rect 397 680 431 682
rect 397 614 431 640
rect 397 606 431 614
rect 397 546 431 566
rect 397 532 431 546
rect 397 478 431 492
rect 397 458 431 478
rect 397 410 431 418
rect 397 384 431 410
rect 241 311 275 342
rect 241 240 275 270
rect 241 236 275 240
rect 320 309 354 343
rect 320 237 354 271
rect 397 342 431 344
rect 397 310 431 342
rect 397 240 431 270
rect 397 236 431 240
rect 553 988 587 1006
rect 553 972 587 988
rect 553 920 587 933
rect 553 899 587 920
rect 553 852 587 860
rect 553 826 587 852
rect 553 784 587 787
rect 553 753 587 784
rect 553 682 587 714
rect 553 680 587 682
rect 553 614 587 640
rect 553 606 587 614
rect 553 546 587 566
rect 553 532 587 546
rect 553 478 587 492
rect 553 458 587 478
rect 553 410 587 418
rect 553 384 587 410
rect 553 342 587 344
rect 553 310 587 342
rect 553 240 587 270
rect 553 236 587 240
rect 709 988 743 1006
rect 709 972 743 988
rect 709 920 743 933
rect 709 899 743 920
rect 709 852 743 860
rect 709 826 743 852
rect 709 784 743 787
rect 709 753 743 784
rect 709 682 743 714
rect 709 680 743 682
rect 709 614 743 640
rect 709 606 743 614
rect 709 546 743 566
rect 709 532 743 546
rect 709 478 743 492
rect 709 458 743 478
rect 709 410 743 418
rect 709 384 743 410
rect 709 342 743 344
rect 709 310 743 342
rect 709 240 743 270
rect 709 236 743 240
rect 865 988 899 1006
rect 865 972 899 988
rect 865 920 899 933
rect 865 899 899 920
rect 865 852 899 860
rect 865 826 899 852
rect 865 784 899 787
rect 865 753 899 784
rect 865 682 899 714
rect 865 680 899 682
rect 865 614 899 640
rect 865 606 899 614
rect 865 546 899 566
rect 865 532 899 546
rect 865 478 899 492
rect 865 458 899 478
rect 865 410 899 418
rect 865 384 899 410
rect 865 342 899 344
rect 865 310 899 342
rect 865 240 899 270
rect 865 236 899 240
rect 1021 1158 1055 1174
rect 1021 1140 1055 1158
rect 1021 1090 1055 1100
rect 1021 1066 1055 1090
rect 1021 1022 1055 1026
rect 1021 992 1055 1022
rect 1021 920 1055 952
rect 1021 918 1055 920
rect 1021 852 1055 878
rect 1021 844 1055 852
rect 1021 784 1055 804
rect 1021 770 1055 784
rect 1021 716 1055 730
rect 1021 696 1055 716
rect 1021 648 1055 656
rect 1021 622 1055 648
rect 1021 580 1055 581
rect 1021 547 1055 580
rect 1021 478 1055 506
rect 1021 472 1055 478
<< metal1 >>
rect 201 1758 1194 1846
rect 201 1724 326 1758
rect 360 1724 402 1758
rect 436 1724 478 1758
rect 512 1724 554 1758
rect 588 1724 630 1758
rect 664 1724 706 1758
rect 740 1724 782 1758
rect 816 1724 858 1758
rect 892 1724 934 1758
rect 968 1724 1011 1758
rect 1045 1724 1194 1758
rect 201 1718 1194 1724
rect 201 1654 247 1718
rect 201 1620 207 1654
rect 241 1620 247 1654
rect 201 1582 247 1620
rect 201 1548 207 1582
rect 241 1548 247 1582
rect 201 1510 247 1548
rect 201 1476 207 1510
rect 241 1476 247 1510
rect 201 1464 247 1476
rect 377 1654 423 1666
rect 377 1620 383 1654
rect 417 1620 423 1654
rect 377 1582 423 1620
rect 377 1548 383 1582
rect 417 1548 423 1582
rect 377 1510 423 1548
rect 377 1476 383 1510
rect 417 1476 423 1510
tri 347 1378 377 1408 se
rect 377 1391 423 1476
rect 553 1654 599 1718
rect 905 1679 951 1718
rect 553 1620 559 1654
rect 593 1620 599 1654
rect 553 1582 599 1620
rect 553 1548 559 1582
rect 593 1548 599 1582
rect 553 1510 599 1548
rect 553 1476 559 1510
rect 593 1476 599 1510
rect 553 1464 599 1476
rect 729 1654 775 1666
rect 729 1620 735 1654
rect 769 1620 775 1654
rect 729 1582 775 1620
rect 729 1548 735 1582
rect 769 1548 775 1582
rect 905 1645 911 1679
rect 945 1645 951 1679
tri 1073 1660 1079 1666 se
rect 1079 1660 1125 1666
tri 1125 1660 1131 1666 sw
rect 905 1597 951 1645
rect 1001 1654 1131 1660
rect 1001 1620 1013 1654
rect 1047 1620 1085 1654
rect 1119 1620 1131 1654
rect 1001 1614 1131 1620
rect 905 1563 911 1597
rect 945 1563 951 1597
rect 905 1551 951 1563
rect 1005 1556 1051 1568
rect 729 1510 775 1548
rect 1005 1522 1011 1556
rect 1045 1522 1051 1556
rect 729 1476 735 1510
rect 769 1476 775 1510
rect 729 1438 775 1476
rect 854 1513 906 1519
rect 854 1449 906 1461
rect 1005 1484 1051 1522
tri 997 1450 1005 1458 se
rect 1005 1450 1011 1484
rect 1045 1450 1051 1484
tri 775 1438 782 1445 sw
rect 729 1435 782 1438
tri 782 1435 785 1438 sw
rect 729 1425 854 1435
tri 729 1415 739 1425 ne
rect 739 1415 854 1425
tri 423 1391 447 1415 sw
tri 739 1391 763 1415 ne
rect 763 1397 854 1415
tri 985 1438 997 1450 se
rect 997 1438 1051 1450
tri 982 1435 985 1438 se
rect 985 1435 1038 1438
rect 906 1425 1038 1435
tri 1038 1425 1051 1438 nw
rect 1079 1565 1131 1614
rect 906 1397 1004 1425
rect 763 1391 1004 1397
tri 1004 1391 1038 1425 nw
tri 1070 1391 1079 1400 se
rect 1079 1391 1125 1565
tri 1125 1559 1131 1565 nw
rect 377 1378 447 1391
rect 142 1362 447 1378
tri 447 1362 476 1391 sw
tri 1041 1362 1070 1391 se
rect 1070 1362 1125 1391
rect 142 1356 1125 1362
rect 142 1333 658 1356
rect 142 1299 154 1333
rect 188 1299 226 1333
rect 260 1322 658 1333
rect 692 1322 748 1356
rect 782 1322 838 1356
rect 872 1322 1125 1356
rect 260 1316 1125 1322
rect 260 1299 273 1316
rect 142 1293 273 1299
tri 273 1293 296 1316 nw
tri 990 1293 1013 1316 ne
rect 1013 1293 1071 1316
tri 1013 1291 1015 1293 ne
rect 1015 1291 1071 1293
tri 1071 1291 1096 1316 nw
rect 1015 1288 1068 1291
tri 1068 1288 1071 1291 nw
tri 252 1232 308 1288 se
rect 308 1282 906 1288
rect 308 1242 854 1282
tri 308 1232 318 1242 nw
tri 213 1193 252 1232 se
rect 252 1193 269 1232
tri 269 1193 308 1232 nw
rect 854 1218 906 1230
tri 201 1181 213 1193 se
rect 213 1181 257 1193
tri 257 1181 269 1193 nw
rect 309 1181 363 1193
tri 196 1176 201 1181 se
rect 201 1176 252 1181
tri 252 1176 257 1181 nw
tri 167 1147 196 1176 se
rect 196 1147 223 1176
tri 223 1147 252 1176 nw
rect 309 1147 320 1181
rect 354 1147 363 1181
rect 854 1160 906 1166
rect 1015 1174 1061 1288
tri 1061 1281 1068 1288 nw
tri 160 1140 167 1147 se
rect 167 1140 216 1147
tri 216 1140 223 1147 nw
tri 152 1132 160 1140 se
rect 160 1132 208 1140
tri 208 1132 216 1140 nw
rect 152 1106 198 1132
tri 198 1122 208 1132 nw
rect 152 1072 158 1106
rect 192 1072 198 1106
rect 309 1109 363 1147
rect 152 1034 198 1072
rect 152 1000 158 1034
rect 192 1000 198 1034
rect 152 988 198 1000
rect 235 1092 281 1104
rect 235 1058 241 1092
rect 275 1058 281 1092
rect 235 1018 281 1058
rect 235 984 241 1018
rect 275 984 281 1018
rect 235 944 281 984
rect 235 910 241 944
rect 275 910 281 944
rect 235 870 281 910
rect 235 836 241 870
rect 275 836 281 870
rect 235 795 281 836
rect 235 761 241 795
rect 275 761 281 795
rect 235 720 281 761
rect 235 710 241 720
rect 152 698 241 710
rect 152 664 158 698
rect 192 686 241 698
rect 275 686 281 720
rect 192 664 281 686
rect 152 645 281 664
rect 152 626 241 645
rect 152 592 158 626
rect 192 611 241 626
rect 275 611 281 645
rect 192 592 281 611
rect 152 580 281 592
rect 235 570 281 580
rect 235 536 241 570
rect 275 536 281 570
rect 235 504 281 536
rect 99 495 281 504
rect 99 492 241 495
rect 99 458 118 492
rect 152 461 241 492
rect 275 461 281 495
rect 152 458 281 461
rect 99 420 281 458
rect 99 414 241 420
rect 99 380 118 414
rect 152 386 241 414
rect 275 386 281 420
rect 152 380 281 386
rect 99 345 281 380
rect 99 336 241 345
rect 99 302 118 336
rect 152 311 241 336
rect 275 311 281 345
rect 152 302 281 311
rect 99 270 281 302
rect 99 258 241 270
rect 99 224 118 258
rect 152 236 241 258
rect 275 236 281 270
rect 152 224 281 236
rect 309 1075 320 1109
rect 354 1075 363 1109
rect 309 343 363 1075
rect 1015 1140 1021 1174
rect 1055 1140 1061 1174
rect 1015 1100 1061 1140
rect 1015 1066 1021 1100
rect 1055 1066 1061 1100
rect 1015 1026 1061 1066
rect 309 309 320 343
rect 354 309 363 343
rect 309 271 363 309
rect 309 237 320 271
rect 354 237 363 271
rect 309 225 363 237
rect 391 1006 437 1018
rect 391 972 397 1006
rect 431 972 437 1006
rect 391 933 437 972
rect 391 899 397 933
rect 431 899 437 933
rect 391 860 437 899
rect 391 826 397 860
rect 431 826 437 860
rect 391 787 437 826
rect 391 753 397 787
rect 431 753 437 787
rect 391 714 437 753
rect 391 680 397 714
rect 431 680 437 714
rect 391 640 437 680
rect 391 606 397 640
rect 431 606 437 640
rect 391 566 437 606
rect 391 532 397 566
rect 431 532 437 566
rect 391 492 437 532
rect 391 458 397 492
rect 431 458 437 492
rect 391 418 437 458
rect 391 384 397 418
rect 431 384 437 418
rect 391 344 437 384
rect 391 310 397 344
rect 431 310 437 344
rect 391 270 437 310
rect 391 236 397 270
rect 431 236 437 270
rect 391 224 437 236
rect 547 1006 593 1018
rect 547 972 553 1006
rect 587 972 593 1006
rect 547 933 593 972
rect 547 899 553 933
rect 587 899 593 933
rect 547 860 593 899
rect 547 826 553 860
rect 587 826 593 860
rect 547 787 593 826
rect 547 753 553 787
rect 587 753 593 787
rect 547 714 593 753
rect 547 680 553 714
rect 587 680 593 714
rect 547 640 593 680
rect 547 606 553 640
rect 587 606 593 640
rect 547 566 593 606
rect 547 532 553 566
rect 587 532 593 566
rect 547 492 593 532
rect 547 458 553 492
rect 587 458 593 492
rect 547 418 593 458
rect 547 384 553 418
rect 587 384 593 418
rect 547 344 593 384
rect 547 310 553 344
rect 587 310 593 344
rect 547 270 593 310
rect 547 236 553 270
rect 587 236 593 270
rect 547 224 593 236
rect 703 1006 749 1018
rect 703 972 709 1006
rect 743 972 749 1006
rect 703 933 749 972
rect 703 899 709 933
rect 743 899 749 933
rect 703 860 749 899
rect 703 826 709 860
rect 743 826 749 860
rect 703 787 749 826
rect 703 753 709 787
rect 743 753 749 787
rect 703 714 749 753
rect 703 680 709 714
rect 743 680 749 714
rect 703 640 749 680
rect 703 606 709 640
rect 743 606 749 640
rect 703 566 749 606
rect 703 532 709 566
rect 743 532 749 566
rect 703 492 749 532
rect 703 458 709 492
rect 743 458 749 492
rect 703 418 749 458
rect 703 384 709 418
rect 743 384 749 418
rect 703 344 749 384
rect 703 310 709 344
rect 743 310 749 344
rect 703 270 749 310
rect 703 236 709 270
rect 743 236 749 270
rect 703 224 749 236
rect 859 1006 905 1018
rect 859 972 865 1006
rect 899 972 905 1006
rect 859 933 905 972
rect 859 899 865 933
rect 899 899 905 933
rect 859 860 905 899
rect 859 826 865 860
rect 899 826 905 860
rect 859 787 905 826
rect 859 753 865 787
rect 899 753 905 787
rect 859 714 905 753
rect 859 680 865 714
rect 899 680 905 714
rect 859 640 905 680
rect 859 606 865 640
rect 899 606 905 640
rect 859 566 905 606
rect 859 532 865 566
rect 899 532 905 566
rect 859 492 905 532
rect 859 458 865 492
rect 899 458 905 492
rect 1015 992 1021 1026
rect 1055 992 1061 1026
rect 1015 952 1061 992
rect 1015 918 1021 952
rect 1055 918 1061 952
rect 1015 878 1061 918
rect 1015 844 1021 878
rect 1055 844 1061 878
rect 1015 804 1061 844
rect 1015 770 1021 804
rect 1055 770 1061 804
rect 1015 730 1061 770
rect 1015 696 1021 730
rect 1055 696 1061 730
rect 1015 656 1061 696
rect 1015 622 1021 656
rect 1055 622 1061 656
rect 1015 581 1061 622
rect 1015 547 1021 581
rect 1055 547 1061 581
rect 1015 506 1061 547
rect 1015 472 1021 506
rect 1055 472 1061 506
rect 1015 460 1061 472
rect 859 418 905 458
rect 859 384 865 418
rect 899 384 905 418
rect 859 344 905 384
rect 859 310 865 344
rect 899 310 905 344
rect 859 270 905 310
rect 859 236 865 270
rect 899 236 905 270
rect 859 224 905 236
rect 99 212 281 224
<< via1 >>
rect 854 1461 906 1513
rect 854 1397 906 1449
rect 854 1230 906 1282
rect 854 1166 906 1218
<< metal2 >>
rect 854 1513 906 1519
rect 854 1449 906 1461
rect 854 1282 906 1397
rect 854 1218 906 1230
rect 854 1160 906 1166
use sky130_fd_pr__nfet_01v8__example_55959141808453  sky130_fd_pr__nfet_01v8__example_55959141808453_0
timestamp 1681267127
transform 1 0 442 0 1 228
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808453  sky130_fd_pr__nfet_01v8__example_55959141808453_1
timestamp 1681267127
transform 1 0 598 0 1 228
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808453  sky130_fd_pr__nfet_01v8__example_55959141808453_2
timestamp 1681267127
transform 1 0 754 0 1 228
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808453  sky130_fd_pr__nfet_01v8__example_55959141808453_3
timestamp 1681267127
transform 1 0 910 0 1 228
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808454  sky130_fd_pr__nfet_01v8__example_55959141808454_0
timestamp 1681267127
transform 1 0 286 0 1 228
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808455  sky130_fd_pr__nfet_01v8__example_55959141808455_0
timestamp 1681267127
transform -1 0 212 0 -1 694
box -19 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808455  sky130_fd_pr__nfet_01v8__example_55959141808455_1
timestamp 1681267127
transform -1 0 212 0 -1 1102
box -19 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808451  sky130_fd_pr__pfet_01v8__example_55959141808451_0
timestamp 1681267127
transform 1 0 974 0 -1 1650
box -19 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808456  sky130_fd_pr__pfet_01v8__example_55959141808456_0
timestamp 1681267127
transform -1 0 900 0 -1 1650
box -1 0 297 1
use sky130_fd_pr__pfet_01v8__example_55959141808457  sky130_fd_pr__pfet_01v8__example_55959141808457_0
timestamp 1681267127
transform 1 0 252 0 -1 1650
box -1 0 297 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_0
timestamp 1681267127
transform 1 0 1013 0 1 1620
box 0 0 1 1
<< labels >>
flabel metal1 s 1049 1323 1077 1351 3 FreeSans 280 180 0 0 OUT
port 1 nsew
flabel metal1 s 485 1739 642 1826 3 FreeSans 520 0 0 0 VPWR
port 2 nsew
flabel metal1 s 157 326 231 434 3 FreeSans 520 0 0 0 VGND
port 3 nsew
flabel locali s 946 109 974 137 3 FreeSans 280 270 0 0 IN1
port 4 nsew
flabel locali s 322 109 350 137 3 FreeSans 280 270 0 0 IN0
port 5 nsew
flabel locali s 634 109 662 137 3 FreeSans 280 270 0 0 IN3
port 6 nsew
flabel locali s 790 109 818 137 3 FreeSans 280 270 0 0 IN2
port 7 nsew
flabel locali s 478 109 506 137 3 FreeSans 280 270 0 0 IN4
port 8 nsew
<< properties >>
string GDS_END 48851806
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 48833828
<< end >>
