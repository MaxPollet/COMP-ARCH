magic
tech sky130A
magscale 1 2
timestamp 1681267127
<< metal4 >>
rect 0 40559 25423 40733
rect 0 40323 287 40559
rect 523 40323 610 40559
rect 846 40323 933 40559
rect 1169 40323 1256 40559
rect 1492 40323 1579 40559
rect 1815 40323 1902 40559
rect 2138 40323 2225 40559
rect 2461 40323 2548 40559
rect 2784 40323 2871 40559
rect 3107 40323 3194 40559
rect 3430 40323 3517 40559
rect 3753 40323 3840 40559
rect 4076 40323 4163 40559
rect 4399 40323 4486 40559
rect 4722 40323 4809 40559
rect 5045 40323 5132 40559
rect 5368 40323 5455 40559
rect 5691 40323 5778 40559
rect 6014 40323 6101 40559
rect 6337 40323 6424 40559
rect 6660 40323 6747 40559
rect 6983 40323 7070 40559
rect 7306 40323 7393 40559
rect 7629 40323 7716 40559
rect 7952 40323 8039 40559
rect 8275 40323 8362 40559
rect 8598 40323 8685 40559
rect 8921 40323 9008 40559
rect 9244 40323 9331 40559
rect 9567 40323 9654 40559
rect 9890 40323 9977 40559
rect 10213 40323 10300 40559
rect 10536 40323 10623 40559
rect 10859 40323 10946 40559
rect 11182 40323 11269 40559
rect 11505 40323 11592 40559
rect 11828 40323 11915 40559
rect 12151 40323 12238 40559
rect 12474 40323 12561 40559
rect 12797 40323 12884 40559
rect 13120 40323 13207 40559
rect 13443 40323 13530 40559
rect 13766 40323 13853 40559
rect 14089 40323 14176 40559
rect 14412 40323 14499 40559
rect 14735 40323 14822 40559
rect 15058 40323 15145 40559
rect 15381 40323 15468 40559
rect 15704 40323 15791 40559
rect 16027 40323 16114 40559
rect 16350 40323 16437 40559
rect 16673 40323 16760 40559
rect 16996 40323 17082 40559
rect 17318 40323 17404 40559
rect 17640 40323 17726 40559
rect 17962 40323 18048 40559
rect 18284 40323 18370 40559
rect 18606 40323 18692 40559
rect 18928 40323 19014 40559
rect 19250 40323 19336 40559
rect 19572 40323 19658 40559
rect 19894 40323 19980 40559
rect 20216 40323 20302 40559
rect 20538 40323 20624 40559
rect 20860 40323 20946 40559
rect 21182 40323 21268 40559
rect 21504 40323 21590 40559
rect 21826 40323 21912 40559
rect 22148 40323 22234 40559
rect 22470 40323 22556 40559
rect 22792 40323 22878 40559
rect 23114 40323 23200 40559
rect 23436 40323 23522 40559
rect 23758 40323 23844 40559
rect 24080 40323 24166 40559
rect 24402 40323 24488 40559
rect 24724 40323 24810 40559
rect 25046 40323 25132 40559
rect 25368 40323 25423 40559
rect 0 40221 25423 40323
rect 0 39985 287 40221
rect 523 39985 610 40221
rect 846 39985 933 40221
rect 1169 39985 1256 40221
rect 1492 39985 1579 40221
rect 1815 39985 1902 40221
rect 2138 39985 2225 40221
rect 2461 39985 2548 40221
rect 2784 39985 2871 40221
rect 3107 39985 3194 40221
rect 3430 39985 3517 40221
rect 3753 39985 3840 40221
rect 4076 39985 4163 40221
rect 4399 39985 4486 40221
rect 4722 39985 4809 40221
rect 5045 39985 5132 40221
rect 5368 39985 5455 40221
rect 5691 39985 5778 40221
rect 6014 39985 6101 40221
rect 6337 39985 6424 40221
rect 6660 39985 6747 40221
rect 6983 39985 7070 40221
rect 7306 39985 7393 40221
rect 7629 39985 7716 40221
rect 7952 39985 8039 40221
rect 8275 39985 8362 40221
rect 8598 39985 8685 40221
rect 8921 39985 9008 40221
rect 9244 39985 9331 40221
rect 9567 39985 9654 40221
rect 9890 39985 9977 40221
rect 10213 39985 10300 40221
rect 10536 39985 10623 40221
rect 10859 39985 10946 40221
rect 11182 39985 11269 40221
rect 11505 39985 11592 40221
rect 11828 39985 11915 40221
rect 12151 39985 12238 40221
rect 12474 39985 12561 40221
rect 12797 39985 12884 40221
rect 13120 39985 13207 40221
rect 13443 39985 13530 40221
rect 13766 39985 13853 40221
rect 14089 39985 14176 40221
rect 14412 39985 14499 40221
rect 14735 39985 14822 40221
rect 15058 39985 15145 40221
rect 15381 39985 15468 40221
rect 15704 39985 15791 40221
rect 16027 39985 16114 40221
rect 16350 39985 16437 40221
rect 16673 39985 16760 40221
rect 16996 39985 17082 40221
rect 17318 39985 17404 40221
rect 17640 39985 17726 40221
rect 17962 39985 18048 40221
rect 18284 39985 18370 40221
rect 18606 39985 18692 40221
rect 18928 39985 19014 40221
rect 19250 39985 19336 40221
rect 19572 39985 19658 40221
rect 19894 39985 19980 40221
rect 20216 39985 20302 40221
rect 20538 39985 20624 40221
rect 20860 39985 20946 40221
rect 21182 39985 21268 40221
rect 21504 39985 21590 40221
rect 21826 39985 21912 40221
rect 22148 39985 22234 40221
rect 22470 39985 22556 40221
rect 22792 39985 22878 40221
rect 23114 39985 23200 40221
rect 23436 39985 23522 40221
rect 23758 39985 23844 40221
rect 24080 39985 24166 40221
rect 24402 39985 24488 40221
rect 24724 39985 24810 40221
rect 25046 39985 25132 40221
rect 25368 39985 25423 40221
rect 0 39900 25423 39985
tri 25423 39900 26256 40733 sw
rect 0 39883 25792 39900
rect 0 39647 287 39883
rect 523 39647 610 39883
rect 846 39647 933 39883
rect 1169 39647 1256 39883
rect 1492 39647 1579 39883
rect 1815 39647 1902 39883
rect 2138 39647 2225 39883
rect 2461 39647 2548 39883
rect 2784 39647 2871 39883
rect 3107 39647 3194 39883
rect 3430 39647 3517 39883
rect 3753 39647 3840 39883
rect 4076 39647 4163 39883
rect 4399 39647 4486 39883
rect 4722 39647 4809 39883
rect 5045 39647 5132 39883
rect 5368 39647 5455 39883
rect 5691 39647 5778 39883
rect 6014 39647 6101 39883
rect 6337 39647 6424 39883
rect 6660 39647 6747 39883
rect 6983 39647 7070 39883
rect 7306 39647 7393 39883
rect 7629 39647 7716 39883
rect 7952 39647 8039 39883
rect 8275 39647 8362 39883
rect 8598 39647 8685 39883
rect 8921 39647 9008 39883
rect 9244 39647 9331 39883
rect 9567 39647 9654 39883
rect 9890 39647 9977 39883
rect 10213 39647 10300 39883
rect 10536 39647 10623 39883
rect 10859 39647 10946 39883
rect 11182 39647 11269 39883
rect 11505 39647 11592 39883
rect 11828 39647 11915 39883
rect 12151 39647 12238 39883
rect 12474 39647 12561 39883
rect 12797 39647 12884 39883
rect 13120 39647 13207 39883
rect 13443 39647 13530 39883
rect 13766 39647 13853 39883
rect 14089 39647 14176 39883
rect 14412 39647 14499 39883
rect 14735 39647 14822 39883
rect 15058 39647 15145 39883
rect 15381 39647 15468 39883
rect 15704 39647 15791 39883
rect 16027 39647 16114 39883
rect 16350 39647 16437 39883
rect 16673 39647 16760 39883
rect 16996 39647 17082 39883
rect 17318 39647 17404 39883
rect 17640 39647 17726 39883
rect 17962 39647 18048 39883
rect 18284 39647 18370 39883
rect 18606 39647 18692 39883
rect 18928 39647 19014 39883
rect 19250 39647 19336 39883
rect 19572 39647 19658 39883
rect 19894 39647 19980 39883
rect 20216 39647 20302 39883
rect 20538 39647 20624 39883
rect 20860 39647 20946 39883
rect 21182 39647 21268 39883
rect 21504 39647 21590 39883
rect 21826 39647 21912 39883
rect 22148 39647 22234 39883
rect 22470 39647 22556 39883
rect 22792 39647 22878 39883
rect 23114 39647 23200 39883
rect 23436 39647 23522 39883
rect 23758 39647 23844 39883
rect 24080 39647 24166 39883
rect 24402 39647 24488 39883
rect 24724 39647 24810 39883
rect 25046 39647 25132 39883
rect 25368 39664 25792 39883
rect 26028 39664 26256 39900
rect 25368 39647 26256 39664
rect 0 39564 26256 39647
rect 0 39545 25792 39564
rect 0 39309 287 39545
rect 523 39309 610 39545
rect 846 39309 933 39545
rect 1169 39309 1256 39545
rect 1492 39309 1579 39545
rect 1815 39309 1902 39545
rect 2138 39309 2225 39545
rect 2461 39309 2548 39545
rect 2784 39309 2871 39545
rect 3107 39309 3194 39545
rect 3430 39309 3517 39545
rect 3753 39309 3840 39545
rect 4076 39309 4163 39545
rect 4399 39309 4486 39545
rect 4722 39309 4809 39545
rect 5045 39309 5132 39545
rect 5368 39309 5455 39545
rect 5691 39309 5778 39545
rect 6014 39309 6101 39545
rect 6337 39309 6424 39545
rect 6660 39309 6747 39545
rect 6983 39309 7070 39545
rect 7306 39309 7393 39545
rect 7629 39309 7716 39545
rect 7952 39309 8039 39545
rect 8275 39309 8362 39545
rect 8598 39309 8685 39545
rect 8921 39309 9008 39545
rect 9244 39309 9331 39545
rect 9567 39309 9654 39545
rect 9890 39309 9977 39545
rect 10213 39309 10300 39545
rect 10536 39309 10623 39545
rect 10859 39309 10946 39545
rect 11182 39309 11269 39545
rect 11505 39309 11592 39545
rect 11828 39309 11915 39545
rect 12151 39309 12238 39545
rect 12474 39309 12561 39545
rect 12797 39309 12884 39545
rect 13120 39309 13207 39545
rect 13443 39309 13530 39545
rect 13766 39309 13853 39545
rect 14089 39309 14176 39545
rect 14412 39309 14499 39545
rect 14735 39309 14822 39545
rect 15058 39309 15145 39545
rect 15381 39309 15468 39545
rect 15704 39309 15791 39545
rect 16027 39309 16114 39545
rect 16350 39309 16437 39545
rect 16673 39309 16760 39545
rect 16996 39309 17082 39545
rect 17318 39309 17404 39545
rect 17640 39309 17726 39545
rect 17962 39309 18048 39545
rect 18284 39309 18370 39545
rect 18606 39309 18692 39545
rect 18928 39309 19014 39545
rect 19250 39309 19336 39545
rect 19572 39309 19658 39545
rect 19894 39309 19980 39545
rect 20216 39309 20302 39545
rect 20538 39309 20624 39545
rect 20860 39309 20946 39545
rect 21182 39309 21268 39545
rect 21504 39309 21590 39545
rect 21826 39309 21912 39545
rect 22148 39309 22234 39545
rect 22470 39309 22556 39545
rect 22792 39309 22878 39545
rect 23114 39309 23200 39545
rect 23436 39309 23522 39545
rect 23758 39309 23844 39545
rect 24080 39309 24166 39545
rect 24402 39309 24488 39545
rect 24724 39309 24810 39545
rect 25046 39309 25132 39545
rect 25368 39328 25792 39545
rect 26028 39328 26256 39564
rect 25368 39309 26256 39328
rect 0 39228 26256 39309
rect 0 39207 25792 39228
rect 0 38971 287 39207
rect 523 38971 610 39207
rect 846 38971 933 39207
rect 1169 38971 1256 39207
rect 1492 38971 1579 39207
rect 1815 38971 1902 39207
rect 2138 38971 2225 39207
rect 2461 38971 2548 39207
rect 2784 38971 2871 39207
rect 3107 38971 3194 39207
rect 3430 38971 3517 39207
rect 3753 38971 3840 39207
rect 4076 38971 4163 39207
rect 4399 38971 4486 39207
rect 4722 38971 4809 39207
rect 5045 38971 5132 39207
rect 5368 38971 5455 39207
rect 5691 38971 5778 39207
rect 6014 38971 6101 39207
rect 6337 38971 6424 39207
rect 6660 38971 6747 39207
rect 6983 38971 7070 39207
rect 7306 38971 7393 39207
rect 7629 38971 7716 39207
rect 7952 38971 8039 39207
rect 8275 38971 8362 39207
rect 8598 38971 8685 39207
rect 8921 38971 9008 39207
rect 9244 38971 9331 39207
rect 9567 38971 9654 39207
rect 9890 38971 9977 39207
rect 10213 38971 10300 39207
rect 10536 38971 10623 39207
rect 10859 38971 10946 39207
rect 11182 38971 11269 39207
rect 11505 38971 11592 39207
rect 11828 38971 11915 39207
rect 12151 38971 12238 39207
rect 12474 38971 12561 39207
rect 12797 38971 12884 39207
rect 13120 38971 13207 39207
rect 13443 38971 13530 39207
rect 13766 38971 13853 39207
rect 14089 38971 14176 39207
rect 14412 38971 14499 39207
rect 14735 38971 14822 39207
rect 15058 38971 15145 39207
rect 15381 38971 15468 39207
rect 15704 38971 15791 39207
rect 16027 38971 16114 39207
rect 16350 38971 16437 39207
rect 16673 38971 16760 39207
rect 16996 38971 17082 39207
rect 17318 38971 17404 39207
rect 17640 38971 17726 39207
rect 17962 38971 18048 39207
rect 18284 38971 18370 39207
rect 18606 38971 18692 39207
rect 18928 38971 19014 39207
rect 19250 38971 19336 39207
rect 19572 38971 19658 39207
rect 19894 38971 19980 39207
rect 20216 38971 20302 39207
rect 20538 38971 20624 39207
rect 20860 38971 20946 39207
rect 21182 38971 21268 39207
rect 21504 38971 21590 39207
rect 21826 38971 21912 39207
rect 22148 38971 22234 39207
rect 22470 38971 22556 39207
rect 22792 38971 22878 39207
rect 23114 38971 23200 39207
rect 23436 38971 23522 39207
rect 23758 38971 23844 39207
rect 24080 38971 24166 39207
rect 24402 38971 24488 39207
rect 24724 38971 24810 39207
rect 25046 38971 25132 39207
rect 25368 38992 25792 39207
rect 26028 38992 26256 39228
rect 25368 38971 26256 38992
rect 0 38961 26256 38971
tri 26256 38961 27195 39900 sw
rect 0 38892 26637 38961
rect 0 38869 25792 38892
rect 0 38633 287 38869
rect 523 38633 610 38869
rect 846 38633 933 38869
rect 1169 38633 1256 38869
rect 1492 38633 1579 38869
rect 1815 38633 1902 38869
rect 2138 38633 2225 38869
rect 2461 38633 2548 38869
rect 2784 38633 2871 38869
rect 3107 38633 3194 38869
rect 3430 38633 3517 38869
rect 3753 38633 3840 38869
rect 4076 38633 4163 38869
rect 4399 38633 4486 38869
rect 4722 38633 4809 38869
rect 5045 38633 5132 38869
rect 5368 38633 5455 38869
rect 5691 38633 5778 38869
rect 6014 38633 6101 38869
rect 6337 38633 6424 38869
rect 6660 38633 6747 38869
rect 6983 38633 7070 38869
rect 7306 38633 7393 38869
rect 7629 38633 7716 38869
rect 7952 38633 8039 38869
rect 8275 38633 8362 38869
rect 8598 38633 8685 38869
rect 8921 38633 9008 38869
rect 9244 38633 9331 38869
rect 9567 38633 9654 38869
rect 9890 38633 9977 38869
rect 10213 38633 10300 38869
rect 10536 38633 10623 38869
rect 10859 38633 10946 38869
rect 11182 38633 11269 38869
rect 11505 38633 11592 38869
rect 11828 38633 11915 38869
rect 12151 38633 12238 38869
rect 12474 38633 12561 38869
rect 12797 38633 12884 38869
rect 13120 38633 13207 38869
rect 13443 38633 13530 38869
rect 13766 38633 13853 38869
rect 14089 38633 14176 38869
rect 14412 38633 14499 38869
rect 14735 38633 14822 38869
rect 15058 38633 15145 38869
rect 15381 38633 15468 38869
rect 15704 38633 15791 38869
rect 16027 38633 16114 38869
rect 16350 38633 16437 38869
rect 16673 38633 16760 38869
rect 16996 38633 17082 38869
rect 17318 38633 17404 38869
rect 17640 38633 17726 38869
rect 17962 38633 18048 38869
rect 18284 38633 18370 38869
rect 18606 38633 18692 38869
rect 18928 38633 19014 38869
rect 19250 38633 19336 38869
rect 19572 38633 19658 38869
rect 19894 38633 19980 38869
rect 20216 38633 20302 38869
rect 20538 38633 20624 38869
rect 20860 38633 20946 38869
rect 21182 38633 21268 38869
rect 21504 38633 21590 38869
rect 21826 38633 21912 38869
rect 22148 38633 22234 38869
rect 22470 38633 22556 38869
rect 22792 38633 22878 38869
rect 23114 38633 23200 38869
rect 23436 38633 23522 38869
rect 23758 38633 23844 38869
rect 24080 38633 24166 38869
rect 24402 38633 24488 38869
rect 24724 38633 24810 38869
rect 25046 38633 25132 38869
rect 25368 38656 25792 38869
rect 26028 38725 26637 38892
rect 26873 38725 27195 38961
rect 26028 38656 27195 38725
rect 25368 38633 27195 38656
rect 0 38625 27195 38633
rect 0 38556 26637 38625
rect 0 38531 25792 38556
rect 0 38295 287 38531
rect 523 38295 610 38531
rect 846 38295 933 38531
rect 1169 38295 1256 38531
rect 1492 38295 1579 38531
rect 1815 38295 1902 38531
rect 2138 38295 2225 38531
rect 2461 38295 2548 38531
rect 2784 38295 2871 38531
rect 3107 38295 3194 38531
rect 3430 38295 3517 38531
rect 3753 38295 3840 38531
rect 4076 38295 4163 38531
rect 4399 38295 4486 38531
rect 4722 38295 4809 38531
rect 5045 38295 5132 38531
rect 5368 38295 5455 38531
rect 5691 38295 5778 38531
rect 6014 38295 6101 38531
rect 6337 38295 6424 38531
rect 6660 38295 6747 38531
rect 6983 38295 7070 38531
rect 7306 38295 7393 38531
rect 7629 38295 7716 38531
rect 7952 38295 8039 38531
rect 8275 38295 8362 38531
rect 8598 38295 8685 38531
rect 8921 38295 9008 38531
rect 9244 38295 9331 38531
rect 9567 38295 9654 38531
rect 9890 38295 9977 38531
rect 10213 38295 10300 38531
rect 10536 38295 10623 38531
rect 10859 38295 10946 38531
rect 11182 38295 11269 38531
rect 11505 38295 11592 38531
rect 11828 38295 11915 38531
rect 12151 38295 12238 38531
rect 12474 38295 12561 38531
rect 12797 38295 12884 38531
rect 13120 38295 13207 38531
rect 13443 38295 13530 38531
rect 13766 38295 13853 38531
rect 14089 38295 14176 38531
rect 14412 38295 14499 38531
rect 14735 38295 14822 38531
rect 15058 38295 15145 38531
rect 15381 38295 15468 38531
rect 15704 38295 15791 38531
rect 16027 38295 16114 38531
rect 16350 38295 16437 38531
rect 16673 38295 16760 38531
rect 16996 38295 17082 38531
rect 17318 38295 17404 38531
rect 17640 38295 17726 38531
rect 17962 38295 18048 38531
rect 18284 38295 18370 38531
rect 18606 38295 18692 38531
rect 18928 38295 19014 38531
rect 19250 38295 19336 38531
rect 19572 38295 19658 38531
rect 19894 38295 19980 38531
rect 20216 38295 20302 38531
rect 20538 38295 20624 38531
rect 20860 38295 20946 38531
rect 21182 38295 21268 38531
rect 21504 38295 21590 38531
rect 21826 38295 21912 38531
rect 22148 38295 22234 38531
rect 22470 38295 22556 38531
rect 22792 38295 22878 38531
rect 23114 38295 23200 38531
rect 23436 38295 23522 38531
rect 23758 38295 23844 38531
rect 24080 38295 24166 38531
rect 24402 38295 24488 38531
rect 24724 38295 24810 38531
rect 25046 38295 25132 38531
rect 25368 38320 25792 38531
rect 26028 38389 26637 38556
rect 26873 38389 27195 38625
rect 26028 38320 27195 38389
rect 25368 38299 27195 38320
tri 27195 38299 27857 38961 sw
rect 25368 38295 27393 38299
rect 0 38289 27393 38295
rect 0 38220 26637 38289
rect 0 38193 25792 38220
rect 0 37957 287 38193
rect 523 37957 610 38193
rect 846 37957 933 38193
rect 1169 37957 1256 38193
rect 1492 37957 1579 38193
rect 1815 37957 1902 38193
rect 2138 37957 2225 38193
rect 2461 37957 2548 38193
rect 2784 37957 2871 38193
rect 3107 37957 3194 38193
rect 3430 37957 3517 38193
rect 3753 37957 3840 38193
rect 4076 37957 4163 38193
rect 4399 37957 4486 38193
rect 4722 37957 4809 38193
rect 5045 37957 5132 38193
rect 5368 37957 5455 38193
rect 5691 37957 5778 38193
rect 6014 37957 6101 38193
rect 6337 37957 6424 38193
rect 6660 37957 6747 38193
rect 6983 37957 7070 38193
rect 7306 37957 7393 38193
rect 7629 37957 7716 38193
rect 7952 37957 8039 38193
rect 8275 37957 8362 38193
rect 8598 37957 8685 38193
rect 8921 37957 9008 38193
rect 9244 37957 9331 38193
rect 9567 37957 9654 38193
rect 9890 37957 9977 38193
rect 10213 37957 10300 38193
rect 10536 37957 10623 38193
rect 10859 37957 10946 38193
rect 11182 37957 11269 38193
rect 11505 37957 11592 38193
rect 11828 37957 11915 38193
rect 12151 37957 12238 38193
rect 12474 37957 12561 38193
rect 12797 37957 12884 38193
rect 13120 37957 13207 38193
rect 13443 37957 13530 38193
rect 13766 37957 13853 38193
rect 14089 37957 14176 38193
rect 14412 37957 14499 38193
rect 14735 37957 14822 38193
rect 15058 37957 15145 38193
rect 15381 37957 15468 38193
rect 15704 37957 15791 38193
rect 16027 37957 16114 38193
rect 16350 37957 16437 38193
rect 16673 37957 16760 38193
rect 16996 37957 17082 38193
rect 17318 37957 17404 38193
rect 17640 37957 17726 38193
rect 17962 37957 18048 38193
rect 18284 37957 18370 38193
rect 18606 37957 18692 38193
rect 18928 37957 19014 38193
rect 19250 37957 19336 38193
rect 19572 37957 19658 38193
rect 19894 37957 19980 38193
rect 20216 37957 20302 38193
rect 20538 37957 20624 38193
rect 20860 37957 20946 38193
rect 21182 37957 21268 38193
rect 21504 37957 21590 38193
rect 21826 37957 21912 38193
rect 22148 37957 22234 38193
rect 22470 37957 22556 38193
rect 22792 37957 22878 38193
rect 23114 37957 23200 38193
rect 23436 37957 23522 38193
rect 23758 37957 23844 38193
rect 24080 37957 24166 38193
rect 24402 37957 24488 38193
rect 24724 37957 24810 38193
rect 25046 37957 25132 38193
rect 25368 37984 25792 38193
rect 26028 38053 26637 38220
rect 26873 38063 27393 38289
rect 27629 38063 27857 38299
rect 26873 38053 27857 38063
rect 26028 37984 27857 38053
rect 25368 37963 27857 37984
rect 25368 37957 27393 37963
rect 0 37953 27393 37957
rect 0 37884 26637 37953
rect 0 37855 25792 37884
rect 0 37619 287 37855
rect 523 37619 610 37855
rect 846 37619 933 37855
rect 1169 37619 1256 37855
rect 1492 37619 1579 37855
rect 1815 37619 1902 37855
rect 2138 37619 2225 37855
rect 2461 37619 2548 37855
rect 2784 37619 2871 37855
rect 3107 37619 3194 37855
rect 3430 37619 3517 37855
rect 3753 37619 3840 37855
rect 4076 37619 4163 37855
rect 4399 37619 4486 37855
rect 4722 37619 4809 37855
rect 5045 37619 5132 37855
rect 5368 37619 5455 37855
rect 5691 37619 5778 37855
rect 6014 37619 6101 37855
rect 6337 37619 6424 37855
rect 6660 37619 6747 37855
rect 6983 37619 7070 37855
rect 7306 37619 7393 37855
rect 7629 37619 7716 37855
rect 7952 37619 8039 37855
rect 8275 37619 8362 37855
rect 8598 37619 8685 37855
rect 8921 37619 9008 37855
rect 9244 37619 9331 37855
rect 9567 37619 9654 37855
rect 9890 37619 9977 37855
rect 10213 37619 10300 37855
rect 10536 37619 10623 37855
rect 10859 37619 10946 37855
rect 11182 37619 11269 37855
rect 11505 37619 11592 37855
rect 11828 37619 11915 37855
rect 12151 37619 12238 37855
rect 12474 37619 12561 37855
rect 12797 37619 12884 37855
rect 13120 37619 13207 37855
rect 13443 37619 13530 37855
rect 13766 37619 13853 37855
rect 14089 37619 14176 37855
rect 14412 37619 14499 37855
rect 14735 37619 14822 37855
rect 15058 37619 15145 37855
rect 15381 37619 15468 37855
rect 15704 37619 15791 37855
rect 16027 37619 16114 37855
rect 16350 37619 16437 37855
rect 16673 37619 16760 37855
rect 16996 37619 17082 37855
rect 17318 37619 17404 37855
rect 17640 37619 17726 37855
rect 17962 37619 18048 37855
rect 18284 37619 18370 37855
rect 18606 37619 18692 37855
rect 18928 37619 19014 37855
rect 19250 37619 19336 37855
rect 19572 37619 19658 37855
rect 19894 37619 19980 37855
rect 20216 37619 20302 37855
rect 20538 37619 20624 37855
rect 20860 37619 20946 37855
rect 21182 37619 21268 37855
rect 21504 37619 21590 37855
rect 21826 37619 21912 37855
rect 22148 37619 22234 37855
rect 22470 37619 22556 37855
rect 22792 37619 22878 37855
rect 23114 37619 23200 37855
rect 23436 37619 23522 37855
rect 23758 37619 23844 37855
rect 24080 37619 24166 37855
rect 24402 37619 24488 37855
rect 24724 37619 24810 37855
rect 25046 37619 25132 37855
rect 25368 37648 25792 37855
rect 26028 37717 26637 37884
rect 26873 37727 27393 37953
rect 27629 37727 27857 37963
rect 26873 37717 27857 37727
rect 26028 37648 27857 37717
rect 25368 37627 27857 37648
rect 25368 37619 27393 37627
rect 0 37617 27393 37619
rect 0 37548 26637 37617
rect 0 37517 25792 37548
rect 0 37281 287 37517
rect 523 37281 610 37517
rect 846 37281 933 37517
rect 1169 37281 1256 37517
rect 1492 37281 1579 37517
rect 1815 37281 1902 37517
rect 2138 37281 2225 37517
rect 2461 37281 2548 37517
rect 2784 37281 2871 37517
rect 3107 37281 3194 37517
rect 3430 37281 3517 37517
rect 3753 37281 3840 37517
rect 4076 37281 4163 37517
rect 4399 37281 4486 37517
rect 4722 37281 4809 37517
rect 5045 37281 5132 37517
rect 5368 37281 5455 37517
rect 5691 37281 5778 37517
rect 6014 37281 6101 37517
rect 6337 37281 6424 37517
rect 6660 37281 6747 37517
rect 6983 37281 7070 37517
rect 7306 37281 7393 37517
rect 7629 37281 7716 37517
rect 7952 37281 8039 37517
rect 8275 37281 8362 37517
rect 8598 37281 8685 37517
rect 8921 37281 9008 37517
rect 9244 37281 9331 37517
rect 9567 37281 9654 37517
rect 9890 37281 9977 37517
rect 10213 37281 10300 37517
rect 10536 37281 10623 37517
rect 10859 37281 10946 37517
rect 11182 37281 11269 37517
rect 11505 37281 11592 37517
rect 11828 37281 11915 37517
rect 12151 37281 12238 37517
rect 12474 37281 12561 37517
rect 12797 37281 12884 37517
rect 13120 37281 13207 37517
rect 13443 37281 13530 37517
rect 13766 37281 13853 37517
rect 14089 37281 14176 37517
rect 14412 37281 14499 37517
rect 14735 37281 14822 37517
rect 15058 37281 15145 37517
rect 15381 37281 15468 37517
rect 15704 37281 15791 37517
rect 16027 37281 16114 37517
rect 16350 37281 16437 37517
rect 16673 37281 16760 37517
rect 16996 37281 17082 37517
rect 17318 37281 17404 37517
rect 17640 37281 17726 37517
rect 17962 37281 18048 37517
rect 18284 37281 18370 37517
rect 18606 37281 18692 37517
rect 18928 37281 19014 37517
rect 19250 37281 19336 37517
rect 19572 37281 19658 37517
rect 19894 37281 19980 37517
rect 20216 37281 20302 37517
rect 20538 37281 20624 37517
rect 20860 37281 20946 37517
rect 21182 37281 21268 37517
rect 21504 37281 21590 37517
rect 21826 37281 21912 37517
rect 22148 37281 22234 37517
rect 22470 37281 22556 37517
rect 22792 37281 22878 37517
rect 23114 37281 23200 37517
rect 23436 37281 23522 37517
rect 23758 37281 23844 37517
rect 24080 37281 24166 37517
rect 24402 37281 24488 37517
rect 24724 37281 24810 37517
rect 25046 37281 25132 37517
rect 25368 37312 25792 37517
rect 26028 37381 26637 37548
rect 26873 37391 27393 37617
rect 27629 37391 27857 37627
rect 26873 37381 27857 37391
rect 26028 37360 27857 37381
tri 27857 37360 28796 38299 sw
rect 26028 37312 28238 37360
rect 25368 37291 28238 37312
rect 25368 37281 27393 37291
rect 0 37211 26637 37281
rect 0 37179 25792 37211
rect 0 36943 287 37179
rect 523 36943 610 37179
rect 846 36943 933 37179
rect 1169 36943 1256 37179
rect 1492 36943 1579 37179
rect 1815 36943 1902 37179
rect 2138 36943 2225 37179
rect 2461 36943 2548 37179
rect 2784 36943 2871 37179
rect 3107 36943 3194 37179
rect 3430 36943 3517 37179
rect 3753 36943 3840 37179
rect 4076 36943 4163 37179
rect 4399 36943 4486 37179
rect 4722 36943 4809 37179
rect 5045 36943 5132 37179
rect 5368 36943 5455 37179
rect 5691 36943 5778 37179
rect 6014 36943 6101 37179
rect 6337 36943 6424 37179
rect 6660 36943 6747 37179
rect 6983 36943 7070 37179
rect 7306 36943 7393 37179
rect 7629 36943 7716 37179
rect 7952 36943 8039 37179
rect 8275 36943 8362 37179
rect 8598 36943 8685 37179
rect 8921 36943 9008 37179
rect 9244 36943 9331 37179
rect 9567 36943 9654 37179
rect 9890 36943 9977 37179
rect 10213 36943 10300 37179
rect 10536 36943 10623 37179
rect 10859 36943 10946 37179
rect 11182 36943 11269 37179
rect 11505 36943 11592 37179
rect 11828 36943 11915 37179
rect 12151 36943 12238 37179
rect 12474 36943 12561 37179
rect 12797 36943 12884 37179
rect 13120 36943 13207 37179
rect 13443 36943 13530 37179
rect 13766 36943 13853 37179
rect 14089 36943 14176 37179
rect 14412 36943 14499 37179
rect 14735 36943 14822 37179
rect 15058 36943 15145 37179
rect 15381 36943 15468 37179
rect 15704 36943 15791 37179
rect 16027 36943 16114 37179
rect 16350 36943 16437 37179
rect 16673 36943 16760 37179
rect 16996 36943 17082 37179
rect 17318 36943 17404 37179
rect 17640 36943 17726 37179
rect 17962 36943 18048 37179
rect 18284 36943 18370 37179
rect 18606 36943 18692 37179
rect 18928 36943 19014 37179
rect 19250 36943 19336 37179
rect 19572 36943 19658 37179
rect 19894 36943 19980 37179
rect 20216 36943 20302 37179
rect 20538 36943 20624 37179
rect 20860 36943 20946 37179
rect 21182 36943 21268 37179
rect 21504 36943 21590 37179
rect 21826 36943 21912 37179
rect 22148 36943 22234 37179
rect 22470 36943 22556 37179
rect 22792 36943 22878 37179
rect 23114 36943 23200 37179
rect 23436 36943 23522 37179
rect 23758 36943 23844 37179
rect 24080 36943 24166 37179
rect 24402 36943 24488 37179
rect 24724 36943 24810 37179
rect 25046 36943 25132 37179
rect 25368 36975 25792 37179
rect 26028 37045 26637 37211
rect 26873 37055 27393 37281
rect 27629 37124 28238 37291
rect 28474 37124 28796 37360
rect 27629 37055 28796 37124
rect 26873 37045 28796 37055
rect 26028 37024 28796 37045
rect 26028 36975 28238 37024
rect 25368 36955 28238 36975
rect 25368 36945 27393 36955
rect 25368 36943 26637 36945
rect 0 36874 26637 36943
rect 0 36841 25792 36874
rect 0 36605 287 36841
rect 523 36605 610 36841
rect 846 36605 933 36841
rect 1169 36605 1256 36841
rect 1492 36605 1579 36841
rect 1815 36605 1902 36841
rect 2138 36605 2225 36841
rect 2461 36605 2548 36841
rect 2784 36605 2871 36841
rect 3107 36605 3194 36841
rect 3430 36605 3517 36841
rect 3753 36605 3840 36841
rect 4076 36605 4163 36841
rect 4399 36605 4486 36841
rect 4722 36605 4809 36841
rect 5045 36605 5132 36841
rect 5368 36605 5455 36841
rect 5691 36605 5778 36841
rect 6014 36605 6101 36841
rect 6337 36605 6424 36841
rect 6660 36605 6747 36841
rect 6983 36605 7070 36841
rect 7306 36605 7393 36841
rect 7629 36605 7716 36841
rect 7952 36605 8039 36841
rect 8275 36605 8362 36841
rect 8598 36605 8685 36841
rect 8921 36605 9008 36841
rect 9244 36605 9331 36841
rect 9567 36605 9654 36841
rect 9890 36605 9977 36841
rect 10213 36605 10300 36841
rect 10536 36605 10623 36841
rect 10859 36605 10946 36841
rect 11182 36605 11269 36841
rect 11505 36605 11592 36841
rect 11828 36605 11915 36841
rect 12151 36605 12238 36841
rect 12474 36605 12561 36841
rect 12797 36605 12884 36841
rect 13120 36605 13207 36841
rect 13443 36605 13530 36841
rect 13766 36605 13853 36841
rect 14089 36605 14176 36841
rect 14412 36605 14499 36841
rect 14735 36605 14822 36841
rect 15058 36605 15145 36841
rect 15381 36605 15468 36841
rect 15704 36605 15791 36841
rect 16027 36605 16114 36841
rect 16350 36605 16437 36841
rect 16673 36605 16760 36841
rect 16996 36605 17082 36841
rect 17318 36605 17404 36841
rect 17640 36605 17726 36841
rect 17962 36605 18048 36841
rect 18284 36605 18370 36841
rect 18606 36605 18692 36841
rect 18928 36605 19014 36841
rect 19250 36605 19336 36841
rect 19572 36605 19658 36841
rect 19894 36605 19980 36841
rect 20216 36605 20302 36841
rect 20538 36605 20624 36841
rect 20860 36605 20946 36841
rect 21182 36605 21268 36841
rect 21504 36605 21590 36841
rect 21826 36605 21912 36841
rect 22148 36605 22234 36841
rect 22470 36605 22556 36841
rect 22792 36605 22878 36841
rect 23114 36605 23200 36841
rect 23436 36605 23522 36841
rect 23758 36605 23844 36841
rect 24080 36605 24166 36841
rect 24402 36605 24488 36841
rect 24724 36605 24810 36841
rect 25046 36605 25132 36841
rect 25368 36638 25792 36841
rect 26028 36709 26637 36874
rect 26873 36719 27393 36945
rect 27629 36788 28238 36955
rect 28474 36788 28796 37024
rect 27629 36719 28796 36788
rect 26873 36709 28796 36719
rect 26028 36698 28796 36709
tri 28796 36698 29458 37360 sw
rect 26028 36688 28994 36698
rect 26028 36638 28238 36688
rect 25368 36619 28238 36638
rect 25368 36609 27393 36619
rect 25368 36605 26637 36609
rect 0 36537 26637 36605
rect 0 36503 25792 36537
rect 0 36267 287 36503
rect 523 36267 610 36503
rect 846 36267 933 36503
rect 1169 36267 1256 36503
rect 1492 36267 1579 36503
rect 1815 36267 1902 36503
rect 2138 36267 2225 36503
rect 2461 36267 2548 36503
rect 2784 36267 2871 36503
rect 3107 36267 3194 36503
rect 3430 36267 3517 36503
rect 3753 36267 3840 36503
rect 4076 36267 4163 36503
rect 4399 36267 4486 36503
rect 4722 36267 4809 36503
rect 5045 36267 5132 36503
rect 5368 36267 5455 36503
rect 5691 36267 5778 36503
rect 6014 36267 6101 36503
rect 6337 36267 6424 36503
rect 6660 36267 6747 36503
rect 6983 36267 7070 36503
rect 7306 36267 7393 36503
rect 7629 36267 7716 36503
rect 7952 36267 8039 36503
rect 8275 36267 8362 36503
rect 8598 36267 8685 36503
rect 8921 36267 9008 36503
rect 9244 36267 9331 36503
rect 9567 36267 9654 36503
rect 9890 36267 9977 36503
rect 10213 36267 10300 36503
rect 10536 36267 10623 36503
rect 10859 36267 10946 36503
rect 11182 36267 11269 36503
rect 11505 36267 11592 36503
rect 11828 36267 11915 36503
rect 12151 36267 12238 36503
rect 12474 36267 12561 36503
rect 12797 36267 12884 36503
rect 13120 36267 13207 36503
rect 13443 36267 13530 36503
rect 13766 36267 13853 36503
rect 14089 36267 14176 36503
rect 14412 36267 14499 36503
rect 14735 36267 14822 36503
rect 15058 36267 15145 36503
rect 15381 36267 15468 36503
rect 15704 36267 15791 36503
rect 16027 36267 16114 36503
rect 16350 36267 16437 36503
rect 16673 36267 16760 36503
rect 16996 36267 17082 36503
rect 17318 36267 17404 36503
rect 17640 36267 17726 36503
rect 17962 36267 18048 36503
rect 18284 36267 18370 36503
rect 18606 36267 18692 36503
rect 18928 36267 19014 36503
rect 19250 36267 19336 36503
rect 19572 36267 19658 36503
rect 19894 36267 19980 36503
rect 20216 36267 20302 36503
rect 20538 36267 20624 36503
rect 20860 36267 20946 36503
rect 21182 36267 21268 36503
rect 21504 36267 21590 36503
rect 21826 36267 21912 36503
rect 22148 36267 22234 36503
rect 22470 36267 22556 36503
rect 22792 36267 22878 36503
rect 23114 36267 23200 36503
rect 23436 36267 23522 36503
rect 23758 36267 23844 36503
rect 24080 36267 24166 36503
rect 24402 36267 24488 36503
rect 24724 36267 24810 36503
rect 25046 36267 25132 36503
rect 25368 36301 25792 36503
rect 26028 36373 26637 36537
rect 26873 36383 27393 36609
rect 27629 36452 28238 36619
rect 28474 36462 28994 36688
rect 29230 36462 29458 36698
rect 28474 36452 29458 36462
rect 27629 36383 29458 36452
rect 26873 36373 29458 36383
rect 26028 36362 29458 36373
rect 26028 36352 28994 36362
rect 26028 36301 28238 36352
rect 25368 36283 28238 36301
rect 25368 36272 27393 36283
rect 25368 36267 26637 36272
rect 0 36200 26637 36267
rect 0 36165 25792 36200
rect 0 35929 287 36165
rect 523 35929 610 36165
rect 846 35929 933 36165
rect 1169 35929 1256 36165
rect 1492 35929 1579 36165
rect 1815 35929 1902 36165
rect 2138 35929 2225 36165
rect 2461 35929 2548 36165
rect 2784 35929 2871 36165
rect 3107 35929 3194 36165
rect 3430 35929 3517 36165
rect 3753 35929 3840 36165
rect 4076 35929 4163 36165
rect 4399 35929 4486 36165
rect 4722 35929 4809 36165
rect 5045 35929 5132 36165
rect 5368 35929 5455 36165
rect 5691 35929 5778 36165
rect 6014 35929 6101 36165
rect 6337 35929 6424 36165
rect 6660 35929 6747 36165
rect 6983 35929 7070 36165
rect 7306 35929 7393 36165
rect 7629 35929 7716 36165
rect 7952 35929 8039 36165
rect 8275 35929 8362 36165
rect 8598 35929 8685 36165
rect 8921 35929 9008 36165
rect 9244 35929 9331 36165
rect 9567 35929 9654 36165
rect 9890 35929 9977 36165
rect 10213 35929 10300 36165
rect 10536 35929 10623 36165
rect 10859 35929 10946 36165
rect 11182 35929 11269 36165
rect 11505 35929 11592 36165
rect 11828 35929 11915 36165
rect 12151 35929 12238 36165
rect 12474 35929 12561 36165
rect 12797 35929 12884 36165
rect 13120 35929 13207 36165
rect 13443 35929 13530 36165
rect 13766 35929 13853 36165
rect 14089 35929 14176 36165
rect 14412 35929 14499 36165
rect 14735 35929 14822 36165
rect 15058 35929 15145 36165
rect 15381 35929 15468 36165
rect 15704 35929 15791 36165
rect 16027 35929 16114 36165
rect 16350 35929 16437 36165
rect 16673 35929 16760 36165
rect 16996 35929 17082 36165
rect 17318 35929 17404 36165
rect 17640 35929 17726 36165
rect 17962 35929 18048 36165
rect 18284 35929 18370 36165
rect 18606 35929 18692 36165
rect 18928 35929 19014 36165
rect 19250 35929 19336 36165
rect 19572 35929 19658 36165
rect 19894 35929 19980 36165
rect 20216 35929 20302 36165
rect 20538 35929 20624 36165
rect 20860 35929 20946 36165
rect 21182 35929 21268 36165
rect 21504 35929 21590 36165
rect 21826 35929 21912 36165
rect 22148 35929 22234 36165
rect 22470 35929 22556 36165
rect 22792 35929 22878 36165
rect 23114 35929 23200 36165
rect 23436 35929 23522 36165
rect 23758 35929 23844 36165
rect 24080 35929 24166 36165
rect 24402 35929 24488 36165
rect 24724 35929 24810 36165
rect 25046 35929 25132 36165
rect 25368 35964 25792 36165
rect 26028 36036 26637 36200
rect 26873 36047 27393 36272
rect 27629 36116 28238 36283
rect 28474 36126 28994 36352
rect 29230 36126 29458 36362
rect 28474 36116 29458 36126
rect 27629 36047 29458 36116
rect 26873 36036 29458 36047
rect 26028 36026 29458 36036
rect 26028 36016 28994 36026
rect 26028 35964 28238 36016
rect 25368 35947 28238 35964
rect 25368 35935 27393 35947
rect 25368 35929 26637 35935
rect 0 35890 26637 35929
tri 23206 33605 25491 35890 ne
rect 25491 35863 26637 35890
rect 25491 35627 25792 35863
rect 26028 35699 26637 35863
rect 26873 35711 27393 35935
rect 27629 35780 28238 35947
rect 28474 35790 28994 36016
rect 29230 35890 29458 36026
tri 29458 35890 30266 36698 sw
rect 29230 35790 30266 35890
rect 28474 35780 30266 35790
rect 27629 35759 30266 35780
rect 27629 35711 29839 35759
rect 26873 35699 29839 35711
rect 26028 35690 29839 35699
rect 26028 35680 28994 35690
rect 26028 35627 28238 35680
rect 25491 35610 28238 35627
rect 25491 35598 27393 35610
rect 25491 35526 26637 35598
rect 25491 35290 25792 35526
rect 26028 35362 26637 35526
rect 26873 35374 27393 35598
rect 27629 35444 28238 35610
rect 28474 35454 28994 35680
rect 29230 35523 29839 35690
rect 30075 35523 30266 35759
rect 29230 35454 30266 35523
rect 28474 35444 30266 35454
rect 27629 35423 30266 35444
rect 27629 35374 29839 35423
rect 26873 35362 29839 35374
rect 26028 35354 29839 35362
rect 26028 35344 28994 35354
rect 26028 35290 28238 35344
rect 25491 35273 28238 35290
rect 25491 35261 27393 35273
rect 25491 35189 26637 35261
rect 25491 34953 25792 35189
rect 26028 35025 26637 35189
rect 26873 35037 27393 35261
rect 27629 35108 28238 35273
rect 28474 35118 28994 35344
rect 29230 35187 29839 35354
rect 30075 35187 30266 35423
rect 29230 35118 30266 35187
rect 28474 35108 30266 35118
rect 27629 35097 30266 35108
tri 30266 35097 31059 35890 sw
rect 27629 35087 30595 35097
rect 27629 35037 29839 35087
rect 26873 35025 29839 35037
rect 26028 35018 29839 35025
rect 26028 35008 28994 35018
rect 26028 34953 28238 35008
rect 25491 34936 28238 34953
rect 25491 34924 27393 34936
rect 25491 34852 26637 34924
rect 25491 34616 25792 34852
rect 26028 34688 26637 34852
rect 26873 34700 27393 34924
rect 27629 34772 28238 34936
rect 28474 34782 28994 35008
rect 29230 34851 29839 35018
rect 30075 34861 30595 35087
rect 30831 34861 31059 35097
rect 30075 34851 31059 34861
rect 29230 34782 31059 34851
rect 28474 34772 31059 34782
rect 27629 34761 31059 34772
rect 27629 34751 30595 34761
rect 27629 34700 29839 34751
rect 26873 34688 29839 34700
rect 26028 34682 29839 34688
rect 26028 34671 28994 34682
rect 26028 34616 28238 34671
rect 25491 34599 28238 34616
rect 25491 34587 27393 34599
rect 25491 34515 26637 34587
rect 25491 34279 25792 34515
rect 26028 34351 26637 34515
rect 26873 34363 27393 34587
rect 27629 34435 28238 34599
rect 28474 34446 28994 34671
rect 29230 34515 29839 34682
rect 30075 34525 30595 34751
rect 30831 34525 31059 34761
rect 30075 34515 31059 34525
rect 29230 34446 31059 34515
rect 28474 34435 31059 34446
rect 27629 34425 31059 34435
rect 27629 34415 30595 34425
rect 27629 34363 29839 34415
rect 26873 34351 29839 34363
rect 26028 34346 29839 34351
rect 26028 34334 28994 34346
rect 26028 34279 28238 34334
rect 25491 34262 28238 34279
rect 25491 34250 27393 34262
rect 25491 34178 26637 34250
rect 25491 33942 25792 34178
rect 26028 34014 26637 34178
rect 26873 34026 27393 34250
rect 27629 34098 28238 34262
rect 28474 34110 28994 34334
rect 29230 34179 29839 34346
rect 30075 34189 30595 34415
rect 30831 34189 31059 34425
rect 30075 34179 31059 34189
rect 29230 34158 31059 34179
tri 31059 34158 31998 35097 sw
rect 29230 34110 31440 34158
rect 28474 34098 31440 34110
rect 27629 34089 31440 34098
rect 27629 34079 30595 34089
rect 27629 34026 29839 34079
rect 26873 34014 29839 34026
rect 26028 34009 29839 34014
rect 26028 33997 28994 34009
rect 26028 33942 28238 33997
rect 25491 33925 28238 33942
rect 25491 33913 27393 33925
rect 25491 33841 26637 33913
rect 25491 33605 25792 33841
rect 26028 33677 26637 33841
rect 26873 33689 27393 33913
rect 27629 33761 28238 33925
rect 28474 33773 28994 33997
rect 29230 33843 29839 34009
rect 30075 33853 30595 34079
rect 30831 33922 31440 34089
rect 31676 33922 31998 34158
rect 30831 33853 31998 33922
rect 30075 33843 31998 33853
rect 29230 33822 31998 33843
rect 29230 33773 31440 33822
rect 28474 33761 31440 33773
rect 27629 33753 31440 33761
rect 27629 33743 30595 33753
rect 27629 33689 29839 33743
rect 26873 33677 29839 33689
rect 26028 33672 29839 33677
rect 26028 33660 28994 33672
rect 26028 33605 28238 33660
tri 25491 32666 26430 33605 ne
rect 26430 33588 28238 33605
rect 26430 33576 27393 33588
rect 26430 33340 26637 33576
rect 26873 33352 27393 33576
rect 27629 33424 28238 33588
rect 28474 33436 28994 33660
rect 29230 33507 29839 33672
rect 30075 33517 30595 33743
rect 30831 33586 31440 33753
rect 31676 33586 31998 33822
rect 30831 33573 31998 33586
tri 31998 33573 32583 34158 sw
rect 30831 33517 32119 33573
rect 30075 33507 32119 33517
rect 29230 33486 32119 33507
rect 29230 33436 31440 33486
rect 28474 33424 31440 33436
rect 27629 33417 31440 33424
rect 27629 33407 30595 33417
rect 27629 33352 29839 33407
rect 26873 33340 29839 33352
rect 26430 33335 29839 33340
rect 26430 33323 28994 33335
rect 26430 33251 28238 33323
rect 26430 33239 27393 33251
rect 26430 33003 26637 33239
rect 26873 33015 27393 33239
rect 27629 33087 28238 33251
rect 28474 33099 28994 33323
rect 29230 33171 29839 33335
rect 30075 33181 30595 33407
rect 30831 33250 31440 33417
rect 31676 33337 32119 33486
rect 32355 33337 32583 33573
rect 31676 33250 32583 33337
rect 30831 33237 32583 33250
rect 30831 33181 32119 33237
rect 30075 33171 32119 33181
rect 29230 33150 32119 33171
rect 29230 33099 31440 33150
rect 28474 33087 31440 33099
rect 27629 33081 31440 33087
rect 27629 33070 30595 33081
rect 27629 33015 29839 33070
rect 26873 33003 29839 33015
rect 26430 32998 29839 33003
rect 26430 32986 28994 32998
rect 26430 32914 28238 32986
rect 26430 32902 27393 32914
rect 26430 32666 26637 32902
rect 26873 32678 27393 32902
rect 27629 32750 28238 32914
rect 28474 32762 28994 32986
rect 29230 32834 29839 32998
rect 30075 32845 30595 33070
rect 30831 32914 31440 33081
rect 31676 33001 32119 33150
rect 32355 33001 32583 33237
rect 31676 32914 32583 33001
rect 30831 32901 32583 32914
rect 30831 32845 32119 32901
rect 30075 32834 32119 32845
rect 29230 32814 32119 32834
rect 29230 32762 31440 32814
rect 28474 32750 31440 32762
rect 27629 32745 31440 32750
rect 27629 32733 30595 32745
rect 27629 32678 29839 32733
rect 26873 32666 29839 32678
tri 26430 32004 27092 32666 ne
rect 27092 32661 29839 32666
rect 27092 32649 28994 32661
rect 27092 32577 28238 32649
rect 27092 32341 27393 32577
rect 27629 32413 28238 32577
rect 28474 32425 28994 32649
rect 29230 32497 29839 32661
rect 30075 32509 30595 32733
rect 30831 32578 31440 32745
rect 31676 32665 32119 32814
rect 32355 32665 32583 32901
rect 31676 32634 32583 32665
tri 32583 32634 33522 33573 sw
rect 31676 32578 32964 32634
rect 30831 32565 32964 32578
rect 30831 32509 32119 32565
rect 30075 32497 32119 32509
rect 29230 32478 32119 32497
rect 29230 32425 31440 32478
rect 28474 32413 31440 32425
rect 27629 32408 31440 32413
rect 27629 32396 30595 32408
rect 27629 32341 29839 32396
rect 27092 32324 29839 32341
rect 27092 32312 28994 32324
rect 27092 32240 28238 32312
rect 27092 32004 27393 32240
rect 27629 32076 28238 32240
rect 28474 32088 28994 32312
rect 29230 32160 29839 32324
rect 30075 32172 30595 32396
rect 30831 32242 31440 32408
rect 31676 32329 32119 32478
rect 32355 32398 32964 32565
rect 33200 32398 33522 32634
rect 32355 32329 33522 32398
rect 31676 32298 33522 32329
rect 31676 32242 32964 32298
rect 30831 32229 32964 32242
rect 30831 32172 32119 32229
rect 30075 32160 32119 32172
rect 29230 32142 32119 32160
rect 29230 32088 31440 32142
rect 28474 32076 31440 32088
rect 27629 32071 31440 32076
rect 27629 32059 30595 32071
rect 27629 32004 29839 32059
tri 27092 31065 28031 32004 ne
rect 28031 31987 29839 32004
rect 28031 31975 28994 31987
rect 28031 31739 28238 31975
rect 28474 31751 28994 31975
rect 29230 31823 29839 31987
rect 30075 31835 30595 32059
rect 30831 31906 31440 32071
rect 31676 31993 32119 32142
rect 32355 32062 32964 32229
rect 33200 32062 33522 32298
rect 32355 31993 33522 32062
rect 31676 31972 33522 31993
tri 33522 31972 34184 32634 sw
rect 31676 31962 33720 31972
rect 31676 31906 32964 31962
rect 30831 31893 32964 31906
rect 30831 31835 32119 31893
rect 30075 31823 32119 31835
rect 29230 31806 32119 31823
rect 29230 31751 31440 31806
rect 28474 31739 31440 31751
rect 28031 31734 31440 31739
rect 28031 31722 30595 31734
rect 28031 31650 29839 31722
rect 28031 31638 28994 31650
rect 28031 31402 28238 31638
rect 28474 31414 28994 31638
rect 29230 31486 29839 31650
rect 30075 31498 30595 31722
rect 30831 31570 31440 31734
rect 31676 31657 32119 31806
rect 32355 31726 32964 31893
rect 33200 31736 33720 31962
rect 33956 31736 34184 31972
rect 33200 31726 34184 31736
rect 32355 31657 34184 31726
rect 31676 31636 34184 31657
rect 31676 31626 33720 31636
rect 31676 31570 32964 31626
rect 30831 31557 32964 31570
rect 30831 31498 32119 31557
rect 30075 31486 32119 31498
rect 29230 31469 32119 31486
rect 29230 31414 31440 31469
rect 28474 31402 31440 31414
rect 28031 31397 31440 31402
rect 28031 31385 30595 31397
rect 28031 31313 29839 31385
rect 28031 31301 28994 31313
rect 28031 31065 28238 31301
rect 28474 31077 28994 31301
rect 29230 31149 29839 31313
rect 30075 31161 30595 31385
rect 30831 31233 31440 31397
rect 31676 31321 32119 31469
rect 32355 31390 32964 31557
rect 33200 31400 33720 31626
rect 33956 31400 34184 31636
rect 33200 31390 34184 31400
rect 32355 31321 34184 31390
rect 31676 31300 34184 31321
rect 31676 31290 33720 31300
rect 31676 31233 32964 31290
rect 30831 31221 32964 31233
rect 30831 31161 32119 31221
rect 30075 31149 32119 31161
rect 29230 31132 32119 31149
rect 29230 31077 31440 31132
rect 28474 31065 31440 31077
tri 28031 30403 28693 31065 ne
rect 28693 31060 31440 31065
rect 28693 31048 30595 31060
rect 28693 30976 29839 31048
rect 28693 30740 28994 30976
rect 29230 30812 29839 30976
rect 30075 30824 30595 31048
rect 30831 30896 31440 31060
rect 31676 30985 32119 31132
rect 32355 31054 32964 31221
rect 33200 31064 33720 31290
rect 33956 31064 34184 31300
rect 33200 31054 34184 31064
rect 32355 31033 34184 31054
tri 34184 31033 35123 31972 sw
rect 32355 30985 34565 31033
rect 31676 30964 34565 30985
rect 31676 30954 33720 30964
rect 31676 30896 32964 30954
rect 30831 30884 32964 30896
rect 30831 30824 32119 30884
rect 30075 30812 32119 30824
rect 29230 30795 32119 30812
rect 29230 30740 31440 30795
rect 28693 30723 31440 30740
rect 28693 30711 30595 30723
rect 28693 30639 29839 30711
rect 28693 30403 28994 30639
rect 29230 30475 29839 30639
rect 30075 30487 30595 30711
rect 30831 30559 31440 30723
rect 31676 30648 32119 30795
rect 32355 30718 32964 30884
rect 33200 30728 33720 30954
rect 33956 30797 34565 30964
rect 34801 30999 35123 31033
tri 35123 30999 35157 31033 sw
rect 34801 30797 35157 30999
rect 33956 30728 35157 30797
rect 33200 30718 35157 30728
rect 32355 30697 35157 30718
rect 32355 30648 34565 30697
rect 31676 30628 34565 30648
rect 31676 30618 33720 30628
rect 31676 30559 32964 30618
rect 30831 30547 32964 30559
rect 30831 30487 32119 30547
rect 30075 30475 32119 30487
rect 29230 30458 32119 30475
rect 29230 30403 31440 30458
tri 28693 29464 29632 30403 ne
rect 29632 30386 31440 30403
rect 29632 30374 30595 30386
rect 29632 30138 29839 30374
rect 30075 30150 30595 30374
rect 30831 30222 31440 30386
rect 31676 30311 32119 30458
rect 32355 30382 32964 30547
rect 33200 30392 33720 30618
rect 33956 30461 34565 30628
rect 34801 30461 35157 30697
rect 33956 30392 35157 30461
rect 33200 30382 35157 30392
rect 32355 30361 35157 30382
rect 32355 30311 34565 30361
rect 31676 30292 34565 30311
rect 31676 30282 33720 30292
rect 31676 30222 32964 30282
rect 30831 30210 32964 30222
rect 30831 30150 32119 30210
rect 30075 30138 32119 30150
rect 29632 30121 32119 30138
rect 29632 30049 31440 30121
rect 29632 30037 30595 30049
rect 29632 29801 29839 30037
rect 30075 29813 30595 30037
rect 30831 29885 31440 30049
rect 31676 29974 32119 30121
rect 32355 30046 32964 30210
rect 33200 30056 33720 30282
rect 33956 30125 34565 30292
rect 34801 30233 35157 30361
tri 35157 30233 35923 30999 sw
rect 34801 30125 35365 30233
rect 33956 30056 35365 30125
rect 33200 30046 35365 30056
rect 32355 30025 35365 30046
rect 32355 29974 34565 30025
rect 31676 29956 34565 29974
rect 31676 29945 33720 29956
rect 31676 29885 32964 29945
rect 30831 29873 32964 29885
rect 30831 29813 32119 29873
rect 30075 29801 32119 29813
rect 29632 29784 32119 29801
rect 29632 29712 31440 29784
rect 29632 29700 30595 29712
rect 29632 29464 29839 29700
rect 30075 29476 30595 29700
rect 30831 29548 31440 29712
rect 31676 29637 32119 29784
rect 32355 29709 32964 29873
rect 33200 29720 33720 29945
rect 33956 29789 34565 29956
rect 34801 29997 35365 30025
rect 35601 29997 35923 30233
rect 34801 29901 35923 29997
rect 34801 29789 35365 29901
rect 33956 29720 35365 29789
rect 33200 29709 35365 29720
rect 32355 29689 35365 29709
rect 32355 29637 34565 29689
rect 31676 29620 34565 29637
rect 31676 29608 33720 29620
rect 31676 29548 32964 29608
rect 30831 29536 32964 29548
rect 30831 29476 32119 29536
rect 30075 29464 32119 29476
tri 29632 28830 30266 29464 ne
rect 30266 29447 32119 29464
rect 30266 29375 31440 29447
rect 30266 29139 30595 29375
rect 30831 29211 31440 29375
rect 31676 29300 32119 29447
rect 32355 29372 32964 29536
rect 33200 29384 33720 29608
rect 33956 29453 34565 29620
rect 34801 29665 35365 29689
rect 35601 29665 35923 29901
rect 34801 29569 35923 29665
rect 34801 29453 35365 29569
rect 33956 29384 35365 29453
rect 33200 29372 35365 29384
rect 32355 29353 35365 29372
rect 32355 29300 34565 29353
rect 31676 29283 34565 29300
rect 31676 29271 33720 29283
rect 31676 29211 32964 29271
rect 30831 29199 32964 29211
rect 30831 29139 32119 29199
rect 30266 29110 32119 29139
rect 30266 29038 31440 29110
rect 30266 28830 30595 29038
tri 30266 28802 30294 28830 ne
rect 30294 28802 30595 28830
rect 30831 28874 31440 29038
rect 31676 28963 32119 29110
rect 32355 29035 32964 29199
rect 33200 29047 33720 29271
rect 33956 29117 34565 29283
rect 34801 29333 35365 29353
rect 35601 29361 35923 29569
tri 35923 29361 36795 30233 sw
rect 35601 29333 36237 29361
rect 34801 29237 36237 29333
rect 34801 29117 35365 29237
rect 33956 29047 35365 29117
rect 33200 29035 35365 29047
rect 32355 29017 35365 29035
rect 32355 28963 34565 29017
rect 31676 28946 34565 28963
rect 31676 28934 33720 28946
rect 31676 28874 32964 28934
rect 30831 28862 32964 28874
rect 30831 28802 32119 28862
tri 30294 27863 31233 28802 ne
rect 31233 28773 32119 28802
rect 31233 28537 31440 28773
rect 31676 28626 32119 28773
rect 32355 28698 32964 28862
rect 33200 28710 33720 28934
rect 33956 28781 34565 28946
rect 34801 29001 35365 29017
rect 35601 29125 36237 29237
rect 36473 29125 36795 29361
rect 35601 29029 36795 29125
rect 35601 29001 36237 29029
rect 34801 28905 36237 29001
rect 34801 28781 35365 28905
rect 33956 28710 35365 28781
rect 33200 28698 35365 28710
rect 32355 28681 35365 28698
rect 32355 28626 34565 28681
rect 31676 28609 34565 28626
rect 31676 28597 33720 28609
rect 31676 28537 32964 28597
rect 31233 28525 32964 28537
rect 31233 28436 32119 28525
rect 31233 28200 31440 28436
rect 31676 28289 32119 28436
rect 32355 28361 32964 28525
rect 33200 28373 33720 28597
rect 33956 28445 34565 28609
rect 34801 28669 35365 28681
rect 35601 28793 36237 28905
rect 36473 28830 36795 29029
tri 36795 28830 37326 29361 sw
rect 36473 28793 37326 28830
rect 35601 28697 37326 28793
rect 35601 28669 36237 28697
rect 34801 28573 36237 28669
rect 34801 28445 35365 28573
rect 33956 28373 35365 28445
rect 33200 28361 35365 28373
rect 32355 28344 35365 28361
rect 32355 28289 34565 28344
rect 31676 28272 34565 28289
rect 31676 28260 33720 28272
rect 31676 28200 32964 28260
rect 31233 28188 32964 28200
rect 31233 28099 32119 28188
rect 31233 27863 31440 28099
rect 31676 27952 32119 28099
rect 32355 28024 32964 28188
rect 33200 28036 33720 28260
rect 33956 28108 34565 28272
rect 34801 28337 35365 28344
rect 35601 28461 36237 28573
rect 36473 28475 37326 28697
tri 37326 28475 37681 28830 sw
rect 36473 28461 37123 28475
rect 35601 28365 37123 28461
rect 35601 28337 36237 28365
rect 34801 28241 36237 28337
rect 34801 28108 35365 28241
rect 33956 28036 35365 28108
rect 33200 28024 35365 28036
rect 32355 28007 35365 28024
rect 32355 27952 34565 28007
rect 31676 27935 34565 27952
rect 31676 27923 33720 27935
rect 31676 27863 32964 27923
tri 31233 27278 31818 27863 ne
rect 31818 27851 32964 27863
rect 31818 27615 32119 27851
rect 32355 27687 32964 27851
rect 33200 27699 33720 27923
rect 33956 27771 34565 27935
rect 34801 28005 35365 28007
rect 35601 28129 36237 28241
rect 36473 28239 37123 28365
rect 37359 28239 37681 28475
rect 36473 28132 37681 28239
rect 36473 28129 37123 28132
rect 35601 28033 37123 28129
rect 35601 28005 36237 28033
rect 34801 27909 36237 28005
rect 34801 27771 35365 27909
rect 33956 27699 35365 27771
rect 33200 27687 35365 27699
rect 32355 27673 35365 27687
rect 35601 27797 36237 27909
rect 36473 27896 37123 28033
rect 37359 27896 37681 28132
rect 36473 27797 37681 27896
rect 35601 27789 37681 27797
rect 35601 27701 37123 27789
rect 35601 27673 36237 27701
rect 32355 27670 36237 27673
rect 32355 27615 34565 27670
rect 31818 27598 34565 27615
rect 31818 27586 33720 27598
rect 31818 27514 32964 27586
rect 31818 27278 32119 27514
rect 32355 27350 32964 27514
rect 33200 27362 33720 27586
rect 33956 27434 34565 27598
rect 34801 27577 36237 27670
rect 34801 27434 35365 27577
rect 33956 27362 35365 27434
rect 33200 27350 35365 27362
rect 32355 27341 35365 27350
rect 35601 27465 36237 27577
rect 36473 27553 37123 27701
rect 37359 27649 37681 27789
tri 37681 27649 38507 28475 sw
rect 37359 27553 37949 27649
rect 36473 27465 37949 27553
rect 35601 27446 37949 27465
rect 35601 27369 37123 27446
rect 35601 27341 36237 27369
rect 32355 27333 36237 27341
rect 32355 27278 34565 27333
tri 31818 26339 32757 27278 ne
rect 32757 27261 34565 27278
rect 32757 27249 33720 27261
rect 32757 27013 32964 27249
rect 33200 27025 33720 27249
rect 33956 27097 34565 27261
rect 34801 27245 36237 27333
rect 34801 27097 35365 27245
rect 33956 27025 35365 27097
rect 33200 27013 35365 27025
rect 32757 27009 35365 27013
rect 35601 27133 36237 27245
rect 36473 27210 37123 27369
rect 37359 27413 37949 27446
rect 38185 27413 38507 27649
rect 37359 27324 38507 27413
rect 37359 27210 37949 27324
rect 36473 27133 37949 27210
rect 35601 27103 37949 27133
rect 35601 27037 37123 27103
rect 35601 27009 36237 27037
rect 32757 26996 36237 27009
rect 32757 26924 34565 26996
rect 32757 26912 33720 26924
rect 32757 26676 32964 26912
rect 33200 26688 33720 26912
rect 33956 26760 34565 26924
rect 34801 26913 36237 26996
rect 34801 26760 35365 26913
rect 33956 26688 35365 26760
rect 33200 26677 35365 26688
rect 35601 26801 36237 26913
rect 36473 26867 37123 27037
rect 37359 27088 37949 27103
rect 38185 27088 38507 27324
rect 37359 26999 38507 27088
rect 37359 26867 37949 26999
rect 36473 26801 37949 26867
rect 35601 26763 37949 26801
rect 38185 26850 38507 26999
tri 38507 26850 39306 27649 sw
rect 38185 26763 38748 26850
rect 35601 26760 38748 26763
rect 35601 26705 37123 26760
rect 35601 26677 36237 26705
rect 33200 26676 36237 26677
rect 32757 26659 36237 26676
rect 32757 26587 34565 26659
rect 32757 26575 33720 26587
rect 32757 26339 32964 26575
rect 33200 26351 33720 26575
rect 33956 26423 34565 26587
rect 34801 26580 36237 26659
rect 34801 26423 35365 26580
rect 33956 26351 35365 26423
rect 33200 26344 35365 26351
rect 35601 26469 36237 26580
rect 36473 26524 37123 26705
rect 37359 26673 38748 26760
rect 37359 26524 37949 26673
rect 36473 26469 37949 26524
rect 35601 26437 37949 26469
rect 38185 26614 38748 26673
rect 38984 26614 39306 26850
rect 38185 26525 39306 26614
rect 38185 26437 38748 26525
rect 35601 26416 38748 26437
rect 35601 26373 37123 26416
rect 35601 26344 36237 26373
rect 33200 26339 36237 26344
tri 32757 25677 33419 26339 ne
rect 33419 26322 36237 26339
rect 33419 26250 34565 26322
rect 33419 26014 33720 26250
rect 33956 26086 34565 26250
rect 34801 26247 36237 26322
rect 34801 26086 35365 26247
rect 33956 26014 35365 26086
rect 33419 26011 35365 26014
rect 35601 26137 36237 26247
rect 36473 26180 37123 26373
rect 37359 26347 38748 26416
rect 37359 26180 37949 26347
rect 36473 26137 37949 26180
rect 35601 26111 37949 26137
rect 38185 26289 38748 26347
rect 38984 26289 39306 26525
rect 38185 26200 39306 26289
rect 38185 26111 38748 26200
rect 35601 26072 38748 26111
rect 35601 26041 37123 26072
rect 35601 26011 36237 26041
rect 33419 25985 36237 26011
rect 33419 25913 34565 25985
rect 33419 25677 33720 25913
rect 33956 25749 34565 25913
rect 34801 25914 36237 25985
rect 34801 25749 35365 25914
rect 33956 25678 35365 25749
rect 35601 25805 36237 25914
rect 36473 25836 37123 26041
rect 37359 26021 38748 26072
rect 37359 25836 37949 26021
rect 36473 25805 37949 25836
rect 35601 25785 37949 25805
rect 38185 25964 38748 26021
rect 38984 26156 39306 26200
tri 39306 26156 40000 26850 sw
rect 38984 25964 40000 26156
rect 38185 25875 40000 25964
rect 38185 25785 38748 25875
rect 35601 25728 38748 25785
rect 35601 25709 37123 25728
rect 35601 25678 36237 25709
rect 33956 25677 36237 25678
tri 33419 24738 34358 25677 ne
rect 34358 25648 36237 25677
rect 34358 25412 34565 25648
rect 34801 25581 36237 25648
rect 34801 25412 35365 25581
rect 34358 25345 35365 25412
rect 35601 25473 36237 25581
rect 36473 25492 37123 25709
rect 37359 25695 38748 25728
rect 37359 25492 37949 25695
rect 36473 25473 37949 25492
rect 35601 25459 37949 25473
rect 38185 25639 38748 25695
rect 38984 25639 40000 25875
rect 38185 25550 40000 25639
rect 38185 25459 38748 25550
rect 35601 25384 38748 25459
rect 35601 25377 37123 25384
rect 35601 25345 36237 25377
rect 34358 25311 36237 25345
rect 34358 25075 34565 25311
rect 34801 25248 36237 25311
rect 34801 25075 35365 25248
rect 34358 25012 35365 25075
rect 35601 25141 36237 25248
rect 36473 25148 37123 25377
rect 37359 25369 38748 25384
rect 37359 25148 37949 25369
rect 36473 25141 37949 25148
rect 35601 25133 37949 25141
rect 38185 25314 38748 25369
rect 38984 25314 40000 25550
rect 38185 25225 40000 25314
rect 38185 25133 38748 25225
rect 35601 25044 38748 25133
rect 35601 25012 36237 25044
rect 34358 24974 36237 25012
rect 34358 24738 34565 24974
rect 34801 24915 36237 24974
rect 34801 24738 35365 24915
tri 34358 23939 35157 24738 ne
rect 35157 24679 35365 24738
rect 35601 24808 36237 24915
rect 36473 25043 38748 25044
rect 36473 25040 37949 25043
rect 36473 24808 37123 25040
rect 35601 24804 37123 24808
rect 37359 24807 37949 25040
rect 38185 24989 38748 25043
rect 38984 24989 40000 25225
rect 38185 24899 40000 24989
rect 38185 24807 38748 24899
rect 37359 24804 38748 24807
rect 35601 24717 38748 24804
rect 35601 24711 37949 24717
rect 35601 24679 36237 24711
rect 35157 24475 36237 24679
rect 36473 24696 37949 24711
rect 36473 24475 37123 24696
rect 35157 24460 37123 24475
rect 37359 24481 37949 24696
rect 38185 24663 38748 24717
rect 38984 24663 40000 24899
rect 38185 24573 40000 24663
rect 38185 24481 38748 24573
rect 37359 24460 38748 24481
rect 35157 24337 38748 24460
rect 38984 24337 40000 24573
rect 35157 23918 40000 24337
rect 35157 23682 35250 23918
rect 35486 23682 35584 23918
rect 35820 23682 35918 23918
rect 36154 23682 36252 23918
rect 36488 23682 36586 23918
rect 36822 23682 36920 23918
rect 37156 23682 37254 23918
rect 37490 23682 37588 23918
rect 37824 23682 37922 23918
rect 38158 23682 38256 23918
rect 38492 23682 38590 23918
rect 38826 23682 38924 23918
rect 39160 23682 39258 23918
rect 39494 23682 39592 23918
rect 39828 23682 40000 23918
rect 35157 23596 40000 23682
rect 35157 23360 35250 23596
rect 35486 23360 35584 23596
rect 35820 23360 35918 23596
rect 36154 23360 36252 23596
rect 36488 23360 36586 23596
rect 36822 23360 36920 23596
rect 37156 23360 37254 23596
rect 37490 23360 37588 23596
rect 37824 23360 37922 23596
rect 38158 23360 38256 23596
rect 38492 23360 38590 23596
rect 38826 23360 38924 23596
rect 39160 23360 39258 23596
rect 39494 23360 39592 23596
rect 39828 23360 40000 23596
rect 35157 23274 40000 23360
rect 35157 23038 35250 23274
rect 35486 23038 35584 23274
rect 35820 23038 35918 23274
rect 36154 23038 36252 23274
rect 36488 23038 36586 23274
rect 36822 23038 36920 23274
rect 37156 23038 37254 23274
rect 37490 23038 37588 23274
rect 37824 23038 37922 23274
rect 38158 23038 38256 23274
rect 38492 23038 38590 23274
rect 38826 23038 38924 23274
rect 39160 23038 39258 23274
rect 39494 23038 39592 23274
rect 39828 23038 40000 23274
rect 35157 22952 40000 23038
rect 35157 22716 35250 22952
rect 35486 22716 35584 22952
rect 35820 22716 35918 22952
rect 36154 22716 36252 22952
rect 36488 22716 36586 22952
rect 36822 22716 36920 22952
rect 37156 22716 37254 22952
rect 37490 22716 37588 22952
rect 37824 22716 37922 22952
rect 38158 22716 38256 22952
rect 38492 22716 38590 22952
rect 38826 22716 38924 22952
rect 39160 22716 39258 22952
rect 39494 22716 39592 22952
rect 39828 22716 40000 22952
rect 35157 22630 40000 22716
rect 35157 22394 35250 22630
rect 35486 22394 35584 22630
rect 35820 22394 35918 22630
rect 36154 22394 36252 22630
rect 36488 22394 36586 22630
rect 36822 22394 36920 22630
rect 37156 22394 37254 22630
rect 37490 22394 37588 22630
rect 37824 22394 37922 22630
rect 38158 22394 38256 22630
rect 38492 22394 38590 22630
rect 38826 22394 38924 22630
rect 39160 22394 39258 22630
rect 39494 22394 39592 22630
rect 39828 22394 40000 22630
rect 35157 22308 40000 22394
rect 35157 22072 35250 22308
rect 35486 22072 35584 22308
rect 35820 22072 35918 22308
rect 36154 22072 36252 22308
rect 36488 22072 36586 22308
rect 36822 22072 36920 22308
rect 37156 22072 37254 22308
rect 37490 22072 37588 22308
rect 37824 22072 37922 22308
rect 38158 22072 38256 22308
rect 38492 22072 38590 22308
rect 38826 22072 38924 22308
rect 39160 22072 39258 22308
rect 39494 22072 39592 22308
rect 39828 22072 40000 22308
rect 35157 21986 40000 22072
rect 35157 21750 35250 21986
rect 35486 21750 35584 21986
rect 35820 21750 35918 21986
rect 36154 21750 36252 21986
rect 36488 21750 36586 21986
rect 36822 21750 36920 21986
rect 37156 21750 37254 21986
rect 37490 21750 37588 21986
rect 37824 21750 37922 21986
rect 38158 21750 38256 21986
rect 38492 21750 38590 21986
rect 38826 21750 38924 21986
rect 39160 21750 39258 21986
rect 39494 21750 39592 21986
rect 39828 21750 40000 21986
rect 35157 21664 40000 21750
rect 35157 21428 35250 21664
rect 35486 21428 35584 21664
rect 35820 21428 35918 21664
rect 36154 21428 36252 21664
rect 36488 21428 36586 21664
rect 36822 21428 36920 21664
rect 37156 21428 37254 21664
rect 37490 21428 37588 21664
rect 37824 21428 37922 21664
rect 38158 21428 38256 21664
rect 38492 21428 38590 21664
rect 38826 21428 38924 21664
rect 39160 21428 39258 21664
rect 39494 21428 39592 21664
rect 39828 21428 40000 21664
rect 35157 21342 40000 21428
rect 35157 21106 35250 21342
rect 35486 21106 35584 21342
rect 35820 21106 35918 21342
rect 36154 21106 36252 21342
rect 36488 21106 36586 21342
rect 36822 21106 36920 21342
rect 37156 21106 37254 21342
rect 37490 21106 37588 21342
rect 37824 21106 37922 21342
rect 38158 21106 38256 21342
rect 38492 21106 38590 21342
rect 38826 21106 38924 21342
rect 39160 21106 39258 21342
rect 39494 21106 39592 21342
rect 39828 21106 40000 21342
rect 35157 21020 40000 21106
rect 35157 20784 35250 21020
rect 35486 20784 35584 21020
rect 35820 20784 35918 21020
rect 36154 20784 36252 21020
rect 36488 20784 36586 21020
rect 36822 20784 36920 21020
rect 37156 20784 37254 21020
rect 37490 20784 37588 21020
rect 37824 20784 37922 21020
rect 38158 20784 38256 21020
rect 38492 20784 38590 21020
rect 38826 20784 38924 21020
rect 39160 20784 39258 21020
rect 39494 20784 39592 21020
rect 39828 20784 40000 21020
rect 35157 20698 40000 20784
rect 35157 20462 35250 20698
rect 35486 20462 35584 20698
rect 35820 20462 35918 20698
rect 36154 20462 36252 20698
rect 36488 20462 36586 20698
rect 36822 20462 36920 20698
rect 37156 20462 37254 20698
rect 37490 20462 37588 20698
rect 37824 20462 37922 20698
rect 38158 20462 38256 20698
rect 38492 20462 38590 20698
rect 38826 20462 38924 20698
rect 39160 20462 39258 20698
rect 39494 20462 39592 20698
rect 39828 20462 40000 20698
rect 35157 20376 40000 20462
rect 35157 20140 35250 20376
rect 35486 20140 35584 20376
rect 35820 20140 35918 20376
rect 36154 20140 36252 20376
rect 36488 20140 36586 20376
rect 36822 20140 36920 20376
rect 37156 20140 37254 20376
rect 37490 20140 37588 20376
rect 37824 20140 37922 20376
rect 38158 20140 38256 20376
rect 38492 20140 38590 20376
rect 38826 20140 38924 20376
rect 39160 20140 39258 20376
rect 39494 20140 39592 20376
rect 39828 20140 40000 20376
rect 35157 20054 40000 20140
rect 35157 19818 35250 20054
rect 35486 19818 35584 20054
rect 35820 19818 35918 20054
rect 36154 19818 36252 20054
rect 36488 19818 36586 20054
rect 36822 19818 36920 20054
rect 37156 19818 37254 20054
rect 37490 19818 37588 20054
rect 37824 19818 37922 20054
rect 38158 19818 38256 20054
rect 38492 19818 38590 20054
rect 38826 19818 38924 20054
rect 39160 19818 39258 20054
rect 39494 19818 39592 20054
rect 39828 19818 40000 20054
rect 0 19536 7764 19733
tri 7764 19536 7961 19733 sw
rect 35157 19732 40000 19818
rect 0 19300 529 19536
rect 765 19300 863 19536
rect 1099 19300 1197 19536
rect 1433 19300 1531 19536
rect 1767 19300 1865 19536
rect 2101 19300 2199 19536
rect 2435 19300 2533 19536
rect 2769 19300 2867 19536
rect 3103 19300 3201 19536
rect 3437 19300 3535 19536
rect 3771 19300 3869 19536
rect 4105 19300 4203 19536
rect 4439 19300 4537 19536
rect 4773 19300 4871 19536
rect 5107 19300 5205 19536
rect 5441 19300 5538 19536
rect 5774 19300 5871 19536
rect 6107 19300 6204 19536
rect 6440 19300 6537 19536
rect 6773 19300 6870 19536
rect 7106 19300 7203 19536
rect 7439 19300 7536 19536
rect 7772 19300 7961 19536
rect 0 19204 7961 19300
rect 0 18968 529 19204
rect 765 18968 863 19204
rect 1099 18968 1197 19204
rect 1433 18968 1531 19204
rect 1767 18968 1865 19204
rect 2101 18968 2199 19204
rect 2435 18968 2533 19204
rect 2769 18968 2867 19204
rect 3103 18968 3201 19204
rect 3437 18968 3535 19204
rect 3771 18968 3869 19204
rect 4105 18968 4203 19204
rect 4439 18968 4537 19204
rect 4773 18968 4871 19204
rect 5107 18968 5205 19204
rect 5441 18968 5538 19204
rect 5774 18968 5871 19204
rect 6107 18968 6204 19204
rect 6440 18968 6537 19204
rect 6773 18968 6870 19204
rect 7106 18968 7203 19204
rect 7439 18968 7536 19204
rect 7772 18968 7961 19204
rect 0 18920 7961 18968
tri 7961 18920 8577 19536 sw
rect 35157 19496 35250 19732
rect 35486 19496 35584 19732
rect 35820 19496 35918 19732
rect 36154 19496 36252 19732
rect 36488 19496 36586 19732
rect 36822 19496 36920 19732
rect 37156 19496 37254 19732
rect 37490 19496 37588 19732
rect 37824 19496 37922 19732
rect 38158 19496 38256 19732
rect 38492 19496 38590 19732
rect 38826 19496 38924 19732
rect 39160 19496 39258 19732
rect 39494 19496 39592 19732
rect 39828 19496 40000 19732
rect 35157 19410 40000 19496
rect 35157 19174 35250 19410
rect 35486 19174 35584 19410
rect 35820 19174 35918 19410
rect 36154 19174 36252 19410
rect 36488 19174 36586 19410
rect 36822 19174 36920 19410
rect 37156 19174 37254 19410
rect 37490 19174 37588 19410
rect 37824 19174 37922 19410
rect 38158 19174 38256 19410
rect 38492 19174 38590 19410
rect 38826 19174 38924 19410
rect 39160 19174 39258 19410
rect 39494 19174 39592 19410
rect 39828 19174 40000 19410
rect 35157 19088 40000 19174
rect 0 18872 8138 18920
rect 0 18636 529 18872
rect 765 18636 863 18872
rect 1099 18636 1197 18872
rect 1433 18636 1531 18872
rect 1767 18636 1865 18872
rect 2101 18636 2199 18872
rect 2435 18636 2533 18872
rect 2769 18636 2867 18872
rect 3103 18636 3201 18872
rect 3437 18636 3535 18872
rect 3771 18636 3869 18872
rect 4105 18636 4203 18872
rect 4439 18636 4537 18872
rect 4773 18636 4871 18872
rect 5107 18636 5205 18872
rect 5441 18636 5538 18872
rect 5774 18636 5871 18872
rect 6107 18636 6204 18872
rect 6440 18636 6537 18872
rect 6773 18636 6870 18872
rect 7106 18636 7203 18872
rect 7439 18636 7536 18872
rect 7772 18684 8138 18872
rect 8374 18684 8577 18920
rect 7772 18636 8577 18684
rect 0 18596 8577 18636
rect 0 18540 8138 18596
rect 0 18304 529 18540
rect 765 18304 863 18540
rect 1099 18304 1197 18540
rect 1433 18304 1531 18540
rect 1767 18304 1865 18540
rect 2101 18304 2199 18540
rect 2435 18304 2533 18540
rect 2769 18304 2867 18540
rect 3103 18304 3201 18540
rect 3437 18304 3535 18540
rect 3771 18304 3869 18540
rect 4105 18304 4203 18540
rect 4439 18304 4537 18540
rect 4773 18304 4871 18540
rect 5107 18304 5205 18540
rect 5441 18304 5538 18540
rect 5774 18304 5871 18540
rect 6107 18304 6204 18540
rect 6440 18304 6537 18540
rect 6773 18304 6870 18540
rect 7106 18304 7203 18540
rect 7439 18304 7536 18540
rect 7772 18360 8138 18540
rect 8374 18360 8577 18596
rect 7772 18304 8577 18360
rect 0 18272 8577 18304
rect 0 18208 8138 18272
rect 0 17972 529 18208
rect 765 17972 863 18208
rect 1099 17972 1197 18208
rect 1433 17972 1531 18208
rect 1767 17972 1865 18208
rect 2101 17972 2199 18208
rect 2435 17972 2533 18208
rect 2769 17972 2867 18208
rect 3103 17972 3201 18208
rect 3437 17972 3535 18208
rect 3771 17972 3869 18208
rect 4105 17972 4203 18208
rect 4439 17972 4537 18208
rect 4773 17972 4871 18208
rect 5107 17972 5205 18208
rect 5441 17972 5538 18208
rect 5774 17972 5871 18208
rect 6107 17972 6204 18208
rect 6440 17972 6537 18208
rect 6773 17972 6870 18208
rect 7106 17972 7203 18208
rect 7439 17972 7536 18208
rect 7772 18036 8138 18208
rect 8374 18223 8577 18272
tri 8577 18223 9274 18920 sw
rect 35157 18852 35250 19088
rect 35486 18852 35584 19088
rect 35820 18852 35918 19088
rect 36154 18852 36252 19088
rect 36488 18852 36586 19088
rect 36822 18852 36920 19088
rect 37156 18852 37254 19088
rect 37490 18852 37588 19088
rect 37824 18852 37922 19088
rect 38158 18852 38256 19088
rect 38492 18852 38590 19088
rect 38826 18852 38924 19088
rect 39160 18852 39258 19088
rect 39494 18852 39592 19088
rect 39828 18852 40000 19088
rect 35157 18766 40000 18852
rect 35157 18530 35250 18766
rect 35486 18530 35584 18766
rect 35820 18530 35918 18766
rect 36154 18530 36252 18766
rect 36488 18530 36586 18766
rect 36822 18530 36920 18766
rect 37156 18530 37254 18766
rect 37490 18530 37588 18766
rect 37824 18530 37922 18766
rect 38158 18530 38256 18766
rect 38492 18530 38590 18766
rect 38826 18530 38924 18766
rect 39160 18530 39258 18766
rect 39494 18530 39592 18766
rect 39828 18530 40000 18766
rect 35157 18444 40000 18530
rect 8374 18036 8835 18223
rect 7772 17987 8835 18036
rect 9071 17987 9274 18223
rect 7772 17972 9274 17987
rect 0 17948 9274 17972
rect 0 17876 8138 17948
rect 0 17640 529 17876
rect 765 17640 863 17876
rect 1099 17640 1197 17876
rect 1433 17640 1531 17876
rect 1767 17640 1865 17876
rect 2101 17640 2199 17876
rect 2435 17640 2533 17876
rect 2769 17640 2867 17876
rect 3103 17640 3201 17876
rect 3437 17640 3535 17876
rect 3771 17640 3869 17876
rect 4105 17640 4203 17876
rect 4439 17640 4537 17876
rect 4773 17640 4871 17876
rect 5107 17640 5205 17876
rect 5441 17640 5538 17876
rect 5774 17640 5871 17876
rect 6107 17640 6204 17876
rect 6440 17640 6537 17876
rect 6773 17640 6870 17876
rect 7106 17640 7203 17876
rect 7439 17640 7536 17876
rect 7772 17712 8138 17876
rect 8374 17899 9274 17948
rect 8374 17712 8835 17899
rect 7772 17663 8835 17712
rect 9071 17663 9274 17899
rect 7772 17640 9274 17663
rect 0 17624 9274 17640
rect 0 17544 8138 17624
rect 0 17308 529 17544
rect 765 17308 863 17544
rect 1099 17308 1197 17544
rect 1433 17308 1531 17544
rect 1767 17308 1865 17544
rect 2101 17308 2199 17544
rect 2435 17308 2533 17544
rect 2769 17308 2867 17544
rect 3103 17308 3201 17544
rect 3437 17308 3535 17544
rect 3771 17308 3869 17544
rect 4105 17308 4203 17544
rect 4439 17308 4537 17544
rect 4773 17308 4871 17544
rect 5107 17308 5205 17544
rect 5441 17308 5538 17544
rect 5774 17308 5871 17544
rect 6107 17308 6204 17544
rect 6440 17308 6537 17544
rect 6773 17308 6870 17544
rect 7106 17308 7203 17544
rect 7439 17308 7536 17544
rect 7772 17388 8138 17544
rect 8374 17575 9274 17624
rect 8374 17388 8835 17575
rect 7772 17339 8835 17388
rect 9071 17564 9274 17575
tri 9274 17564 9933 18223 sw
rect 35157 18208 35250 18444
rect 35486 18208 35584 18444
rect 35820 18208 35918 18444
rect 36154 18208 36252 18444
rect 36488 18208 36586 18444
rect 36822 18208 36920 18444
rect 37156 18208 37254 18444
rect 37490 18208 37588 18444
rect 37824 18208 37922 18444
rect 38158 18208 38256 18444
rect 38492 18208 38590 18444
rect 38826 18208 38924 18444
rect 39160 18208 39258 18444
rect 39494 18208 39592 18444
rect 39828 18208 40000 18444
rect 35157 18122 40000 18208
rect 35157 17886 35250 18122
rect 35486 17886 35584 18122
rect 35820 17886 35918 18122
rect 36154 17886 36252 18122
rect 36488 17886 36586 18122
rect 36822 17886 36920 18122
rect 37156 17886 37254 18122
rect 37490 17886 37588 18122
rect 37824 17886 37922 18122
rect 38158 17886 38256 18122
rect 38492 17886 38590 18122
rect 38826 17886 38924 18122
rect 39160 17886 39258 18122
rect 39494 17886 39592 18122
rect 39828 17886 40000 18122
rect 35157 17800 40000 17886
rect 35157 17564 35250 17800
rect 35486 17564 35584 17800
rect 35820 17564 35918 17800
rect 36154 17564 36252 17800
rect 36488 17564 36586 17800
rect 36822 17564 36920 17800
rect 37156 17564 37254 17800
rect 37490 17564 37588 17800
rect 37824 17564 37922 17800
rect 38158 17564 38256 17800
rect 38492 17564 38590 17800
rect 38826 17564 38924 17800
rect 39160 17564 39258 17800
rect 39494 17564 39592 17800
rect 39828 17564 40000 17800
rect 9071 17339 9494 17564
rect 7772 17328 9494 17339
rect 9730 17328 9933 17564
rect 7772 17308 9933 17328
rect 0 17300 9933 17308
rect 0 17212 8138 17300
rect 0 16976 529 17212
rect 765 16976 863 17212
rect 1099 16976 1197 17212
rect 1433 16976 1531 17212
rect 1767 16976 1865 17212
rect 2101 16976 2199 17212
rect 2435 16976 2533 17212
rect 2769 16976 2867 17212
rect 3103 16976 3201 17212
rect 3437 16976 3535 17212
rect 3771 16976 3869 17212
rect 4105 16976 4203 17212
rect 4439 16976 4537 17212
rect 4773 16976 4871 17212
rect 5107 16976 5205 17212
rect 5441 16976 5538 17212
rect 5774 16976 5871 17212
rect 6107 16976 6204 17212
rect 6440 16976 6537 17212
rect 6773 16976 6870 17212
rect 7106 16976 7203 17212
rect 7439 16976 7536 17212
rect 7772 17064 8138 17212
rect 8374 17251 9933 17300
rect 8374 17064 8835 17251
rect 7772 17015 8835 17064
rect 9071 17240 9933 17251
rect 9071 17015 9494 17240
rect 7772 17004 9494 17015
rect 9730 17004 9933 17240
rect 7772 16976 9933 17004
rect 0 16880 8138 16976
rect 0 16644 529 16880
rect 765 16644 863 16880
rect 1099 16644 1197 16880
rect 1433 16644 1531 16880
rect 1767 16644 1865 16880
rect 2101 16644 2199 16880
rect 2435 16644 2533 16880
rect 2769 16644 2867 16880
rect 3103 16644 3201 16880
rect 3437 16644 3535 16880
rect 3771 16644 3869 16880
rect 4105 16644 4203 16880
rect 4439 16644 4537 16880
rect 4773 16644 4871 16880
rect 5107 16644 5205 16880
rect 5441 16644 5538 16880
rect 5774 16644 5871 16880
rect 6107 16644 6204 16880
rect 6440 16644 6537 16880
rect 6773 16644 6870 16880
rect 7106 16644 7203 16880
rect 7439 16644 7536 16880
rect 7772 16740 8138 16880
rect 8374 16927 9933 16976
rect 8374 16740 8835 16927
rect 7772 16691 8835 16740
rect 9071 16916 9933 16927
rect 9071 16691 9494 16916
rect 7772 16680 9494 16691
rect 9730 16867 9933 16916
tri 9933 16867 10630 17564 sw
rect 35157 17478 40000 17564
rect 35157 17242 35250 17478
rect 35486 17242 35584 17478
rect 35820 17242 35918 17478
rect 36154 17242 36252 17478
rect 36488 17242 36586 17478
rect 36822 17242 36920 17478
rect 37156 17242 37254 17478
rect 37490 17242 37588 17478
rect 37824 17242 37922 17478
rect 38158 17242 38256 17478
rect 38492 17242 38590 17478
rect 38826 17242 38924 17478
rect 39160 17242 39258 17478
rect 39494 17242 39592 17478
rect 39828 17242 40000 17478
rect 35157 17156 40000 17242
rect 35157 16920 35250 17156
rect 35486 16920 35584 17156
rect 35820 16920 35918 17156
rect 36154 16920 36252 17156
rect 36488 16920 36586 17156
rect 36822 16920 36920 17156
rect 37156 16920 37254 17156
rect 37490 16920 37588 17156
rect 37824 16920 37922 17156
rect 38158 16920 38256 17156
rect 38492 16920 38590 17156
rect 38826 16920 38924 17156
rect 39160 16920 39258 17156
rect 39494 16920 39592 17156
rect 39828 16920 40000 17156
rect 9730 16680 10191 16867
rect 7772 16652 10191 16680
rect 7772 16644 8138 16652
rect 0 16548 8138 16644
rect 0 16312 529 16548
rect 765 16312 863 16548
rect 1099 16312 1197 16548
rect 1433 16312 1531 16548
rect 1767 16312 1865 16548
rect 2101 16312 2199 16548
rect 2435 16312 2533 16548
rect 2769 16312 2867 16548
rect 3103 16312 3201 16548
rect 3437 16312 3535 16548
rect 3771 16312 3869 16548
rect 4105 16312 4203 16548
rect 4439 16312 4537 16548
rect 4773 16312 4871 16548
rect 5107 16312 5205 16548
rect 5441 16312 5538 16548
rect 5774 16312 5871 16548
rect 6107 16312 6204 16548
rect 6440 16312 6537 16548
rect 6773 16312 6870 16548
rect 7106 16312 7203 16548
rect 7439 16312 7536 16548
rect 7772 16416 8138 16548
rect 8374 16631 10191 16652
rect 10427 16631 10630 16867
rect 8374 16603 10630 16631
rect 8374 16416 8835 16603
rect 7772 16367 8835 16416
rect 9071 16592 10630 16603
rect 9071 16367 9494 16592
rect 7772 16356 9494 16367
rect 9730 16543 10630 16592
rect 9730 16356 10191 16543
rect 7772 16328 10191 16356
rect 7772 16312 8138 16328
rect 0 16216 8138 16312
rect 0 15980 529 16216
rect 765 15980 863 16216
rect 1099 15980 1197 16216
rect 1433 15980 1531 16216
rect 1767 15980 1865 16216
rect 2101 15980 2199 16216
rect 2435 15980 2533 16216
rect 2769 15980 2867 16216
rect 3103 15980 3201 16216
rect 3437 15980 3535 16216
rect 3771 15980 3869 16216
rect 4105 15980 4203 16216
rect 4439 15980 4537 16216
rect 4773 15980 4871 16216
rect 5107 15980 5205 16216
rect 5441 15980 5538 16216
rect 5774 15980 5871 16216
rect 6107 15980 6204 16216
rect 6440 15980 6537 16216
rect 6773 15980 6870 16216
rect 7106 15980 7203 16216
rect 7439 15980 7536 16216
rect 7772 16092 8138 16216
rect 8374 16307 10191 16328
rect 10427 16307 10630 16543
rect 8374 16279 10630 16307
rect 8374 16092 8835 16279
rect 7772 16043 8835 16092
rect 9071 16268 10630 16279
rect 9071 16043 9494 16268
rect 7772 16032 9494 16043
rect 9730 16219 10630 16268
rect 9730 16032 10191 16219
rect 7772 16004 10191 16032
rect 7772 15980 8138 16004
rect 0 15884 8138 15980
rect 0 15648 529 15884
rect 765 15648 863 15884
rect 1099 15648 1197 15884
rect 1433 15648 1531 15884
rect 1767 15648 1865 15884
rect 2101 15648 2199 15884
rect 2435 15648 2533 15884
rect 2769 15648 2867 15884
rect 3103 15648 3201 15884
rect 3437 15648 3535 15884
rect 3771 15648 3869 15884
rect 4105 15648 4203 15884
rect 4439 15648 4537 15884
rect 4773 15648 4871 15884
rect 5107 15648 5205 15884
rect 5441 15648 5538 15884
rect 5774 15648 5871 15884
rect 6107 15648 6204 15884
rect 6440 15648 6537 15884
rect 6773 15648 6870 15884
rect 7106 15648 7203 15884
rect 7439 15648 7536 15884
rect 7772 15768 8138 15884
rect 8374 15983 10191 16004
rect 10427 16188 10630 16219
tri 10630 16188 11309 16867 sw
rect 35157 16834 40000 16920
rect 35157 16598 35250 16834
rect 35486 16598 35584 16834
rect 35820 16598 35918 16834
rect 36154 16598 36252 16834
rect 36488 16598 36586 16834
rect 36822 16598 36920 16834
rect 37156 16598 37254 16834
rect 37490 16598 37588 16834
rect 37824 16598 37922 16834
rect 38158 16598 38256 16834
rect 38492 16598 38590 16834
rect 38826 16598 38924 16834
rect 39160 16598 39258 16834
rect 39494 16598 39592 16834
rect 39828 16598 40000 16834
rect 35157 16512 40000 16598
rect 35157 16276 35250 16512
rect 35486 16276 35584 16512
rect 35820 16276 35918 16512
rect 36154 16276 36252 16512
rect 36488 16276 36586 16512
rect 36822 16276 36920 16512
rect 37156 16276 37254 16512
rect 37490 16276 37588 16512
rect 37824 16276 37922 16512
rect 38158 16276 38256 16512
rect 38492 16276 38590 16512
rect 38826 16276 38924 16512
rect 39160 16276 39258 16512
rect 39494 16276 39592 16512
rect 39828 16276 40000 16512
rect 35157 16190 40000 16276
rect 10427 15983 10870 16188
rect 8374 15955 10870 15983
rect 8374 15768 8835 15955
rect 7772 15719 8835 15768
rect 9071 15952 10870 15955
rect 11106 15952 11309 16188
rect 9071 15944 11309 15952
rect 9071 15719 9494 15944
rect 7772 15708 9494 15719
rect 9730 15895 11309 15944
rect 9730 15708 10191 15895
rect 7772 15680 10191 15708
rect 7772 15648 8138 15680
rect 0 15552 8138 15648
rect 0 15316 529 15552
rect 765 15316 863 15552
rect 1099 15316 1197 15552
rect 1433 15316 1531 15552
rect 1767 15316 1865 15552
rect 2101 15316 2199 15552
rect 2435 15316 2533 15552
rect 2769 15316 2867 15552
rect 3103 15316 3201 15552
rect 3437 15316 3535 15552
rect 3771 15316 3869 15552
rect 4105 15316 4203 15552
rect 4439 15316 4537 15552
rect 4773 15316 4871 15552
rect 5107 15316 5205 15552
rect 5441 15316 5538 15552
rect 5774 15316 5871 15552
rect 6107 15316 6204 15552
rect 6440 15316 6537 15552
rect 6773 15316 6870 15552
rect 7106 15316 7203 15552
rect 7439 15316 7536 15552
rect 7772 15444 8138 15552
rect 8374 15659 10191 15680
rect 10427 15864 11309 15895
rect 10427 15659 10870 15864
rect 8374 15631 10870 15659
rect 8374 15444 8835 15631
rect 7772 15395 8835 15444
rect 9071 15628 10870 15631
rect 11106 15628 11309 15864
rect 9071 15620 11309 15628
rect 9071 15395 9494 15620
rect 7772 15384 9494 15395
rect 9730 15571 11309 15620
rect 9730 15384 10191 15571
rect 7772 15356 10191 15384
rect 7772 15316 8138 15356
rect 0 15220 8138 15316
rect 0 14984 529 15220
rect 765 14984 863 15220
rect 1099 14984 1197 15220
rect 1433 14984 1531 15220
rect 1767 14984 1865 15220
rect 2101 14984 2199 15220
rect 2435 14984 2533 15220
rect 2769 14984 2867 15220
rect 3103 14984 3201 15220
rect 3437 14984 3535 15220
rect 3771 14984 3869 15220
rect 4105 14984 4203 15220
rect 4439 14984 4537 15220
rect 4773 14984 4871 15220
rect 5107 14984 5205 15220
rect 5441 14984 5538 15220
rect 5774 14984 5871 15220
rect 6107 14984 6204 15220
rect 6440 14984 6537 15220
rect 6773 14984 6870 15220
rect 7106 14984 7203 15220
rect 7439 14984 7536 15220
rect 7772 15120 8138 15220
rect 8374 15335 10191 15356
rect 10427 15555 11309 15571
tri 11309 15555 11942 16188 sw
rect 35157 15954 35250 16190
rect 35486 15954 35584 16190
rect 35820 15954 35918 16190
rect 36154 15954 36252 16190
rect 36488 15954 36586 16190
rect 36822 15954 36920 16190
rect 37156 15954 37254 16190
rect 37490 15954 37588 16190
rect 37824 15954 37922 16190
rect 38158 15954 38256 16190
rect 38492 15954 38590 16190
rect 38826 15954 38924 16190
rect 39160 15954 39258 16190
rect 39494 15954 39592 16190
rect 39828 15954 40000 16190
rect 35157 15868 40000 15954
rect 35157 15632 35250 15868
rect 35486 15632 35584 15868
rect 35820 15632 35918 15868
rect 36154 15632 36252 15868
rect 36488 15632 36586 15868
rect 36822 15632 36920 15868
rect 37156 15632 37254 15868
rect 37490 15632 37588 15868
rect 37824 15632 37922 15868
rect 38158 15632 38256 15868
rect 38492 15632 38590 15868
rect 38826 15632 38924 15868
rect 39160 15632 39258 15868
rect 39494 15632 39592 15868
rect 39828 15632 40000 15868
rect 10427 15540 11942 15555
rect 10427 15335 10870 15540
rect 8374 15307 10870 15335
rect 8374 15120 8835 15307
rect 7772 15071 8835 15120
rect 9071 15304 10870 15307
rect 11106 15491 11942 15540
rect 11106 15304 11567 15491
rect 9071 15296 11567 15304
rect 9071 15071 9494 15296
rect 7772 15060 9494 15071
rect 9730 15255 11567 15296
rect 11803 15255 11942 15491
rect 9730 15247 11942 15255
rect 9730 15060 10191 15247
rect 7772 15032 10191 15060
rect 7772 14984 8138 15032
rect 0 14796 8138 14984
rect 8374 15011 10191 15032
rect 10427 15216 11942 15247
rect 10427 15011 10870 15216
rect 8374 14983 10870 15011
rect 8374 14796 8835 14983
rect 0 14747 8835 14796
rect 9071 14980 10870 14983
rect 11106 15167 11942 15216
rect 11106 14980 11567 15167
rect 9071 14972 11567 14980
rect 9071 14747 9494 14972
rect 0 14740 9494 14747
tri 5699 14440 5999 14740 ne
rect 5999 14736 9494 14740
rect 9730 14931 11567 14972
rect 11803 14931 11942 15167
rect 9730 14923 11942 14931
rect 9730 14736 10191 14923
rect 5999 14708 10191 14736
rect 5999 14472 8138 14708
rect 8374 14687 10191 14708
rect 10427 14892 11942 14923
rect 10427 14687 10870 14892
rect 8374 14659 10870 14687
rect 8374 14472 8835 14659
rect 5999 14440 8835 14472
rect 0 14390 5612 14440
rect 0 14154 296 14390
rect 532 14154 627 14390
rect 863 14154 958 14390
rect 1194 14154 1289 14390
rect 1525 14154 1620 14390
rect 1856 14154 1951 14390
rect 2187 14154 2282 14390
rect 2518 14154 2613 14390
rect 2849 14154 2944 14390
rect 3180 14154 3275 14390
rect 3511 14154 3606 14390
rect 3842 14154 3936 14390
rect 4172 14154 4266 14390
rect 4502 14154 4596 14390
rect 4832 14154 4926 14390
rect 5162 14154 5256 14390
rect 5492 14154 5612 14390
rect 0 14092 5612 14154
tri 5612 14092 5960 14440 sw
tri 5999 14092 6347 14440 ne
rect 6347 14423 8835 14440
rect 9071 14656 10870 14659
rect 11106 14843 11942 14892
rect 11106 14656 11567 14843
rect 9071 14648 11567 14656
rect 9071 14423 9494 14648
rect 6347 14412 9494 14423
rect 9730 14607 11567 14648
rect 11803 14832 11942 14843
tri 11942 14832 12665 15555 sw
rect 35157 15546 40000 15632
rect 35157 15310 35250 15546
rect 35486 15310 35584 15546
rect 35820 15310 35918 15546
rect 36154 15310 36252 15546
rect 36488 15310 36586 15546
rect 36822 15310 36920 15546
rect 37156 15310 37254 15546
rect 37490 15310 37588 15546
rect 37824 15310 37922 15546
rect 38158 15310 38256 15546
rect 38492 15310 38590 15546
rect 38826 15310 38924 15546
rect 39160 15310 39258 15546
rect 39494 15310 39592 15546
rect 39828 15310 40000 15546
rect 35157 15224 40000 15310
rect 35157 14988 35250 15224
rect 35486 14988 35584 15224
rect 35820 14988 35918 15224
rect 36154 14988 36252 15224
rect 36488 14988 36586 15224
rect 36822 14988 36920 15224
rect 37156 14988 37254 15224
rect 37490 14988 37588 15224
rect 37824 14988 37922 15224
rect 38158 14988 38256 15224
rect 38492 14988 38590 15224
rect 38826 14988 38924 15224
rect 39160 14988 39258 15224
rect 39494 14988 39592 15224
rect 39828 14988 40000 15224
rect 35157 14902 40000 14988
rect 11803 14607 12226 14832
rect 9730 14599 12226 14607
rect 9730 14412 10191 14599
rect 6347 14384 10191 14412
rect 6347 14148 8138 14384
rect 8374 14363 10191 14384
rect 10427 14596 12226 14599
rect 12462 14596 12665 14832
rect 10427 14568 12665 14596
rect 10427 14363 10870 14568
rect 8374 14335 10870 14363
rect 8374 14148 8835 14335
rect 6347 14099 8835 14148
rect 9071 14332 10870 14335
rect 11106 14519 12665 14568
rect 11106 14332 11567 14519
rect 9071 14324 11567 14332
rect 9071 14099 9494 14324
rect 6347 14092 9494 14099
rect 0 13856 5581 14092
rect 5817 14053 5960 14092
tri 5960 14053 5999 14092 sw
tri 6347 14053 6386 14092 ne
rect 6386 14088 9494 14092
rect 9730 14283 11567 14324
rect 11803 14508 12665 14519
rect 11803 14283 12226 14508
rect 9730 14275 12226 14283
rect 9730 14088 10191 14275
rect 6386 14060 10191 14088
rect 6386 14053 8138 14060
rect 5817 13937 5999 14053
tri 5999 13937 6115 14053 sw
tri 6386 13937 6502 14053 ne
rect 6502 13937 8138 14053
rect 5817 13856 6115 13937
rect 0 13836 6115 13856
rect 0 13600 296 13836
rect 532 13600 627 13836
rect 863 13600 958 13836
rect 1194 13600 1289 13836
rect 1525 13600 1620 13836
rect 1856 13600 1951 13836
rect 2187 13600 2282 13836
rect 2518 13600 2613 13836
rect 2849 13600 2944 13836
rect 3180 13600 3275 13836
rect 3511 13600 3606 13836
rect 3842 13600 3936 13836
rect 4172 13600 4266 13836
rect 4502 13600 4596 13836
rect 4832 13600 4926 13836
rect 5162 13600 5256 13836
rect 5492 13688 6115 13836
tri 6115 13688 6364 13937 sw
tri 6502 13688 6751 13937 ne
rect 6751 13824 8138 13937
rect 8374 14039 10191 14060
rect 10427 14272 12226 14275
rect 12462 14272 12665 14508
rect 10427 14244 12665 14272
rect 10427 14039 10870 14244
rect 8374 14011 10870 14039
rect 8374 13824 8835 14011
rect 6751 13775 8835 13824
rect 9071 14008 10870 14011
rect 11106 14195 12665 14244
rect 11106 14008 11567 14195
rect 9071 14000 11567 14008
rect 9071 13775 9494 14000
rect 6751 13764 9494 13775
rect 9730 13959 11567 14000
rect 11803 14184 12665 14195
rect 11803 13959 12226 14184
rect 9730 13951 12226 13959
rect 9730 13764 10191 13951
rect 6751 13736 10191 13764
rect 6751 13688 8138 13736
rect 5492 13600 5985 13688
rect 0 13550 5985 13600
tri 5241 13270 5521 13550 ne
rect 5521 13545 5985 13550
rect 5521 13309 5581 13545
rect 5817 13452 5985 13545
rect 6221 13550 6364 13688
tri 6364 13550 6502 13688 sw
tri 6751 13550 6889 13688 ne
rect 6889 13550 8138 13688
rect 6221 13452 6502 13550
rect 5817 13309 6502 13452
rect 5521 13282 6502 13309
tri 6502 13282 6770 13550 sw
tri 6889 13282 7157 13550 ne
rect 7157 13500 8138 13550
rect 8374 13715 10191 13736
rect 10427 13948 12226 13951
rect 12462 14135 12665 14184
tri 12665 14135 13362 14832 sw
rect 35157 14666 35250 14902
rect 35486 14666 35584 14902
rect 35820 14666 35918 14902
rect 36154 14666 36252 14902
rect 36488 14666 36586 14902
rect 36822 14666 36920 14902
rect 37156 14666 37254 14902
rect 37490 14666 37588 14902
rect 37824 14666 37922 14902
rect 38158 14666 38256 14902
rect 38492 14666 38590 14902
rect 38826 14666 38924 14902
rect 39160 14666 39258 14902
rect 39494 14666 39592 14902
rect 39828 14666 40000 14902
rect 35157 14580 40000 14666
rect 35157 14344 35250 14580
rect 35486 14344 35584 14580
rect 35820 14344 35918 14580
rect 36154 14344 36252 14580
rect 36488 14344 36586 14580
rect 36822 14344 36920 14580
rect 37156 14344 37254 14580
rect 37490 14344 37588 14580
rect 37824 14344 37922 14580
rect 38158 14344 38256 14580
rect 38492 14344 38590 14580
rect 38826 14344 38924 14580
rect 39160 14344 39258 14580
rect 39494 14344 39592 14580
rect 39828 14344 40000 14580
rect 35157 14258 40000 14344
rect 12462 13948 12923 14135
rect 10427 13920 12923 13948
rect 10427 13715 10870 13920
rect 8374 13687 10870 13715
rect 8374 13500 8835 13687
rect 7157 13451 8835 13500
rect 9071 13684 10870 13687
rect 11106 13899 12923 13920
rect 13159 13899 13362 14135
rect 11106 13871 13362 13899
rect 11106 13684 11567 13871
rect 9071 13676 11567 13684
rect 9071 13451 9494 13676
rect 7157 13440 9494 13451
rect 9730 13635 11567 13676
rect 11803 13860 13362 13871
rect 11803 13635 12226 13860
rect 9730 13627 12226 13635
rect 9730 13440 10191 13627
rect 7157 13412 10191 13440
rect 7157 13282 8138 13412
rect 5521 13270 6391 13282
rect 0 13215 5133 13270
rect 0 12979 325 13215
rect 561 12979 830 13215
rect 1066 12979 1335 13215
rect 1571 12979 1840 13215
rect 2076 12979 2345 13215
rect 2581 12979 2850 13215
rect 3086 12979 3354 13215
rect 3590 12979 3858 13215
rect 4094 12979 4362 13215
rect 4598 12979 4866 13215
rect 5102 12979 5133 13215
rect 0 12882 5133 12979
tri 5133 12882 5521 13270 sw
tri 5521 12882 5909 13270 ne
rect 5909 13141 6391 13270
rect 5909 12905 5985 13141
rect 6221 13046 6391 13141
rect 6627 13163 6770 13282
tri 6770 13163 6889 13282 sw
tri 7157 13163 7276 13282 ne
rect 7276 13176 8138 13282
rect 8374 13391 10191 13412
rect 10427 13624 12226 13627
rect 12462 13811 13362 13860
rect 12462 13624 12923 13811
rect 10427 13596 12923 13624
rect 10427 13391 10870 13596
rect 8374 13363 10870 13391
rect 8374 13176 8835 13363
rect 7276 13163 8835 13176
rect 6627 13063 6889 13163
tri 6889 13063 6989 13163 sw
tri 7276 13063 7376 13163 ne
rect 7376 13127 8835 13163
rect 9071 13360 10870 13363
rect 11106 13575 12923 13596
rect 13159 13575 13362 13811
rect 11106 13547 13362 13575
rect 11106 13360 11567 13547
rect 9071 13352 11567 13360
rect 9071 13127 9494 13352
rect 7376 13116 9494 13127
rect 9730 13311 11567 13352
rect 11803 13536 13362 13547
rect 11803 13311 12226 13536
rect 9730 13303 12226 13311
rect 9730 13116 10191 13303
rect 7376 13088 10191 13116
rect 7376 13063 8138 13088
rect 6627 13046 6989 13063
rect 6221 12905 6989 13046
rect 5909 12882 6989 12905
rect 0 12842 5521 12882
rect 0 12677 5220 12842
rect 0 12441 325 12677
rect 561 12441 830 12677
rect 1066 12441 1335 12677
rect 1571 12441 1840 12677
rect 2076 12441 2345 12677
rect 2581 12441 2850 12677
rect 3086 12441 3354 12677
rect 3590 12441 3858 12677
rect 4094 12441 4362 12677
rect 4598 12441 4866 12677
rect 5102 12606 5220 12677
rect 5456 12606 5521 12842
rect 5102 12564 5521 12606
tri 5521 12564 5839 12882 sw
tri 5909 12564 6227 12882 ne
rect 6227 12878 6989 12882
tri 6989 12878 7174 13063 sw
tri 7376 12878 7561 13063 ne
rect 7561 12878 8138 13063
rect 6227 12735 6795 12878
rect 6227 12564 6391 12735
rect 5102 12478 5839 12564
rect 5102 12441 5581 12478
rect 0 12380 5581 12441
tri 4761 12176 4965 12380 ne
rect 4965 12295 5581 12380
rect 4965 12176 5220 12295
tri 4965 12080 5061 12176 ne
rect 5061 12080 5220 12176
rect 0 12014 4635 12080
tri 4635 12014 4701 12080 sw
tri 5061 12014 5127 12080 ne
rect 5127 12059 5220 12080
rect 5456 12242 5581 12295
rect 5817 12289 5839 12478
tri 5839 12289 6114 12564 sw
tri 6227 12499 6292 12564 ne
rect 6292 12499 6391 12564
rect 6627 12642 6795 12735
rect 7031 12676 7174 12878
tri 7174 12676 7376 12878 sw
tri 7561 12676 7763 12878 ne
rect 7763 12852 8138 12878
rect 8374 13067 10191 13088
rect 10427 13300 12226 13303
rect 12462 13511 13362 13536
tri 13362 13511 13986 14135 sw
rect 35157 14022 35250 14258
rect 35486 14022 35584 14258
rect 35820 14022 35918 14258
rect 36154 14022 36252 14258
rect 36488 14022 36586 14258
rect 36822 14022 36920 14258
rect 37156 14022 37254 14258
rect 37490 14022 37588 14258
rect 37824 14022 37922 14258
rect 38158 14022 38256 14258
rect 38492 14022 38590 14258
rect 38826 14022 38924 14258
rect 39160 14022 39258 14258
rect 39494 14022 39592 14258
rect 39828 14022 40000 14258
rect 35157 13936 40000 14022
rect 35157 13700 35250 13936
rect 35486 13700 35584 13936
rect 35820 13700 35918 13936
rect 36154 13700 36252 13936
rect 36488 13700 36586 13936
rect 36822 13700 36920 13936
rect 37156 13700 37254 13936
rect 37490 13700 37588 13936
rect 37824 13700 37922 13936
rect 38158 13700 38256 13936
rect 38492 13700 38590 13936
rect 38826 13700 38924 13936
rect 39160 13700 39258 13936
rect 39494 13700 39592 13936
rect 39828 13700 40000 13936
rect 35157 13614 40000 13700
rect 12462 13487 13547 13511
rect 12462 13300 12923 13487
rect 10427 13272 12923 13300
rect 10427 13067 10870 13272
rect 8374 13039 10870 13067
rect 8374 12852 8835 13039
rect 7763 12803 8835 12852
rect 9071 13036 10870 13039
rect 11106 13251 12923 13272
rect 13159 13275 13547 13487
rect 13783 13275 13986 13511
rect 13159 13251 13986 13275
rect 11106 13223 13986 13251
rect 11106 13036 11567 13223
rect 9071 13028 11567 13036
rect 9071 12803 9494 13028
rect 7763 12792 9494 12803
rect 9730 12987 11567 13028
rect 11803 13212 13986 13223
rect 11803 12987 12226 13212
rect 9730 12979 12226 12987
rect 9730 12792 10191 12979
rect 7763 12763 10191 12792
rect 7763 12676 8138 12763
rect 7031 12642 7376 12676
rect 6627 12499 7376 12642
tri 6292 12289 6502 12499 ne
rect 6502 12479 7376 12499
tri 7376 12479 7573 12676 sw
tri 7763 12527 7912 12676 ne
rect 7912 12527 8138 12676
rect 8374 12743 10191 12763
rect 10427 12976 12226 12979
rect 12462 13187 13986 13212
rect 12462 13163 13547 13187
rect 12462 12976 12923 13163
rect 10427 12948 12923 12976
rect 10427 12743 10870 12948
rect 8374 12715 10870 12743
rect 8374 12527 8835 12715
tri 7912 12479 7960 12527 ne
rect 7960 12479 8835 12527
rect 9071 12712 10870 12715
rect 11106 12927 12923 12948
rect 13159 12951 13547 13163
rect 13783 12951 13986 13187
rect 13159 12927 13986 12951
rect 11106 12899 13986 12927
rect 11106 12712 11567 12899
rect 9071 12704 11567 12712
rect 9071 12479 9494 12704
rect 6502 12331 7194 12479
rect 6502 12289 6795 12331
rect 5817 12242 6114 12289
rect 5456 12176 6114 12242
tri 6114 12176 6227 12289 sw
tri 6502 12176 6615 12289 ne
rect 6615 12176 6795 12289
rect 5456 12074 6227 12176
rect 5456 12059 5985 12074
rect 5127 12014 5985 12059
tri 4607 12008 4613 12014 ne
rect 4613 12008 4701 12014
tri 4701 12008 4707 12014 sw
tri 5127 12008 5133 12014 ne
rect 5133 12008 5985 12014
tri 4613 11954 4667 12008 ne
rect 4667 11954 4707 12008
tri 4707 11954 4761 12008 sw
tri 5133 11954 5187 12008 ne
rect 5187 11954 5985 12008
rect 0 11920 4582 11954
tri 4582 11920 4616 11954 sw
tri 4667 11920 4701 11954 ne
rect 4701 11920 4761 11954
tri 4761 11920 4795 11954 sw
tri 5187 11920 5221 11954 ne
rect 5221 11931 5985 11954
rect 5221 11920 5581 11931
rect 0 11835 4616 11920
tri 4616 11835 4701 11920 sw
tri 4701 11835 4786 11920 ne
rect 4786 11835 4795 11920
rect 0 11826 4701 11835
tri 4701 11826 4710 11835 sw
tri 4786 11826 4795 11835 ne
tri 4795 11826 4889 11920 sw
tri 5221 11826 5315 11920 ne
rect 5315 11826 5581 11920
rect 0 11741 4710 11826
tri 4710 11741 4795 11826 sw
tri 4795 11741 4880 11826 ne
rect 4880 11741 4889 11826
rect 0 11732 4795 11741
tri 4795 11732 4804 11741 sw
tri 4880 11732 4889 11741 ne
tri 4889 11732 4983 11826 sw
tri 5315 11814 5327 11826 ne
rect 5327 11814 5581 11826
tri 5327 11732 5409 11814 ne
rect 5409 11732 5581 11814
rect 0 11647 4804 11732
tri 4804 11647 4889 11732 sw
tri 4889 11647 4974 11732 ne
rect 4974 11647 4983 11732
rect 0 11638 4889 11647
tri 4889 11638 4898 11647 sw
tri 4974 11638 4983 11647 ne
tri 4983 11638 5077 11732 sw
tri 5409 11638 5503 11732 ne
rect 5503 11695 5581 11732
rect 5817 11838 5985 11931
rect 6221 11838 6227 12074
rect 5817 11788 6227 11838
tri 6227 11788 6615 12176 sw
tri 6615 12095 6696 12176 ne
rect 6696 12095 6795 12176
rect 7031 12243 7194 12331
rect 7430 12289 7573 12479
tri 7573 12289 7763 12479 sw
tri 7960 12289 8150 12479 ne
rect 8150 12468 9494 12479
rect 9730 12663 11567 12704
rect 11803 12888 13986 12899
rect 11803 12663 12226 12888
rect 9730 12655 12226 12663
rect 9730 12468 10191 12655
rect 8150 12419 10191 12468
rect 10427 12652 12226 12655
rect 12462 12863 13986 12888
rect 12462 12839 13547 12863
rect 12462 12652 12923 12839
rect 10427 12624 12923 12652
rect 10427 12419 10870 12624
rect 8150 12391 10870 12419
rect 8150 12289 8835 12391
rect 7430 12243 7763 12289
rect 7031 12095 7763 12243
tri 6696 11788 7003 12095 ne
rect 7003 12075 7763 12095
tri 7763 12075 7977 12289 sw
tri 8150 12075 8364 12289 ne
rect 8364 12155 8835 12289
rect 9071 12388 10870 12391
rect 11106 12603 12923 12624
rect 13159 12627 13547 12839
rect 13783 12814 13986 12863
tri 13986 12814 14683 13511 sw
rect 35157 13378 35250 13614
rect 35486 13378 35584 13614
rect 35820 13378 35918 13614
rect 36154 13378 36252 13614
rect 36488 13378 36586 13614
rect 36822 13378 36920 13614
rect 37156 13378 37254 13614
rect 37490 13378 37588 13614
rect 37824 13378 37922 13614
rect 38158 13378 38256 13614
rect 38492 13378 38590 13614
rect 38826 13378 38924 13614
rect 39160 13378 39258 13614
rect 39494 13378 39592 13614
rect 39828 13378 40000 13614
rect 35157 13292 40000 13378
rect 35157 13056 35250 13292
rect 35486 13056 35584 13292
rect 35820 13056 35918 13292
rect 36154 13056 36252 13292
rect 36488 13056 36586 13292
rect 36822 13056 36920 13292
rect 37156 13056 37254 13292
rect 37490 13056 37588 13292
rect 37824 13056 37922 13292
rect 38158 13056 38256 13292
rect 38492 13056 38590 13292
rect 38826 13056 38924 13292
rect 39160 13056 39258 13292
rect 39494 13056 39592 13292
rect 39828 13056 40000 13292
rect 35157 12970 40000 13056
rect 13783 12627 14244 12814
rect 13159 12603 14244 12627
rect 11106 12578 14244 12603
rect 14480 12578 14683 12814
rect 11106 12575 14683 12578
rect 11106 12388 11567 12575
rect 9071 12380 11567 12388
rect 9071 12155 9494 12380
rect 8364 12144 9494 12155
rect 9730 12339 11567 12380
rect 11803 12564 14683 12575
rect 11803 12339 12226 12564
rect 9730 12331 12226 12339
rect 9730 12144 10191 12331
rect 8364 12095 10191 12144
rect 10427 12328 12226 12331
rect 12462 12539 14683 12564
rect 12462 12515 13547 12539
rect 12462 12328 12923 12515
rect 10427 12300 12923 12328
rect 10427 12095 10870 12300
rect 8364 12075 10870 12095
rect 7003 11932 7598 12075
rect 7003 11788 7194 11932
rect 5817 11695 6615 11788
rect 5503 11690 6615 11695
tri 6615 11690 6713 11788 sw
tri 7003 11690 7101 11788 ne
rect 7101 11696 7194 11788
rect 7430 11839 7598 11932
rect 7834 11902 7977 12075
tri 7977 11902 8150 12075 sw
tri 8364 11902 8537 12075 ne
rect 8537 12066 10870 12075
rect 8537 11902 8835 12066
rect 7834 11839 8150 11902
rect 7430 11802 8150 11839
tri 8150 11802 8250 11902 sw
tri 8537 11802 8637 11902 ne
rect 8637 11830 8835 11902
rect 9071 12064 10870 12066
rect 11106 12279 12923 12300
rect 13159 12303 13547 12515
rect 13783 12492 14683 12539
rect 13783 12303 14244 12492
rect 13159 12279 14244 12303
rect 11106 12256 14244 12279
rect 14480 12256 14683 12492
rect 11106 12251 14683 12256
rect 11106 12064 11567 12251
rect 9071 12056 11567 12064
rect 9071 11830 9494 12056
rect 8637 11820 9494 11830
rect 9730 12015 11567 12056
rect 11803 12240 14683 12251
rect 11803 12015 12226 12240
rect 9730 12007 12226 12015
rect 9730 11820 10191 12007
rect 8637 11802 10191 11820
rect 7430 11696 8250 11802
rect 7101 11690 8250 11696
rect 5503 11668 6713 11690
rect 5503 11638 6391 11668
rect 0 11553 4898 11638
tri 4898 11553 4983 11638 sw
tri 4983 11553 5068 11638 ne
rect 5068 11553 5077 11638
rect 0 11544 4983 11553
tri 4983 11544 4992 11553 sw
tri 5068 11544 5077 11553 ne
tri 5077 11544 5171 11638 sw
tri 5503 11544 5597 11638 ne
rect 5597 11544 6391 11638
rect 0 11459 4992 11544
tri 4992 11459 5077 11544 sw
tri 5077 11459 5162 11544 ne
rect 5162 11459 5171 11544
rect 0 11450 5077 11459
tri 5077 11450 5086 11459 sw
tri 5162 11450 5171 11459 ne
tri 5171 11450 5265 11544 sw
tri 5597 11450 5691 11544 ne
rect 5691 11527 6391 11544
rect 5691 11450 5985 11527
rect 0 11365 5086 11450
tri 5086 11365 5171 11450 sw
tri 5171 11365 5256 11450 ne
rect 5256 11388 5265 11450
tri 5265 11388 5327 11450 sw
tri 5691 11388 5753 11450 ne
rect 5753 11388 5985 11450
rect 5256 11365 5327 11388
rect 0 11358 5171 11365
tri 4336 11298 4396 11358 ne
rect 4396 11356 5171 11358
tri 5171 11356 5180 11365 sw
tri 5256 11356 5265 11365 ne
rect 5265 11356 5327 11365
tri 5327 11356 5359 11388 sw
tri 5753 11356 5785 11388 ne
rect 5785 11356 5985 11388
rect 4396 11298 5180 11356
rect 0 11212 4310 11298
tri 4310 11212 4396 11298 sw
tri 4396 11212 4482 11298 ne
rect 4482 11294 5180 11298
tri 5180 11294 5242 11356 sw
tri 5265 11294 5327 11356 ne
rect 5327 11294 5359 11356
rect 4482 11262 5242 11294
tri 5242 11262 5274 11294 sw
tri 5327 11262 5359 11294 ne
tri 5359 11262 5453 11356 sw
tri 5785 11262 5879 11356 ne
rect 5879 11291 5985 11356
rect 6221 11432 6391 11527
rect 6627 11432 6713 11668
rect 6221 11302 6713 11432
tri 6713 11302 7101 11690 sw
tri 7101 11302 7489 11690 ne
rect 7489 11664 8250 11690
rect 7489 11528 8009 11664
rect 7489 11302 7598 11528
rect 6221 11291 7101 11302
rect 5879 11262 7101 11291
rect 4482 11212 5274 11262
rect 0 11209 4396 11212
tri 4396 11209 4399 11212 sw
tri 4482 11209 4485 11212 ne
rect 4485 11209 5274 11212
tri 5274 11209 5327 11262 sw
tri 5359 11209 5412 11262 ne
rect 5412 11209 5453 11262
tri 5453 11209 5506 11262 sw
tri 5879 11209 5932 11262 ne
rect 5932 11209 6800 11262
rect 0 11148 4399 11209
tri 4399 11148 4460 11209 sw
tri 4485 11148 4546 11209 ne
rect 4546 11168 5327 11209
tri 5327 11168 5368 11209 sw
tri 5412 11168 5453 11209 ne
rect 5453 11168 5506 11209
tri 5506 11168 5547 11209 sw
tri 5932 11168 5973 11209 ne
rect 5973 11168 6800 11209
rect 4546 11148 5368 11168
rect 0 11112 4460 11148
tri 4460 11112 4496 11148 sw
tri 4546 11112 4582 11148 ne
rect 4582 11112 5368 11148
rect 0 11062 4496 11112
tri 4496 11062 4546 11112 sw
tri 4582 11062 4632 11112 ne
rect 4632 11083 5368 11112
tri 5368 11083 5453 11168 sw
tri 5453 11083 5538 11168 ne
rect 5538 11083 5547 11168
rect 4632 11074 5453 11083
tri 5453 11074 5462 11083 sw
tri 5538 11074 5547 11083 ne
tri 5547 11074 5641 11168 sw
tri 5973 11074 6067 11168 ne
rect 6067 11121 6800 11168
rect 6067 11074 6391 11121
rect 4632 11062 5462 11074
tri 4212 11002 4272 11062 ne
rect 4272 11002 4546 11062
rect 0 10977 4187 11002
tri 4187 10977 4212 11002 sw
tri 4272 10977 4297 11002 ne
rect 4297 10977 4546 11002
rect 0 10906 4212 10977
tri 4212 10906 4283 10977 sw
tri 4297 10906 4368 10977 ne
rect 4368 10976 4546 10977
tri 4546 10976 4632 11062 sw
tri 4632 10976 4718 11062 ne
rect 4718 10989 5462 11062
tri 5462 10989 5547 11074 sw
tri 5547 10989 5632 11074 ne
rect 5632 10989 5641 11074
rect 4718 10980 5547 10989
tri 5547 10980 5556 10989 sw
tri 5632 10980 5641 10989 ne
tri 5641 10980 5735 11074 sw
tri 6067 10980 6161 11074 ne
rect 6161 10980 6391 11074
rect 4718 10976 5556 10980
rect 4368 10907 4632 10976
tri 4632 10907 4701 10976 sw
tri 4718 10907 4787 10976 ne
rect 4787 10914 5556 10976
tri 5556 10914 5622 10980 sw
tri 5641 10914 5707 10980 ne
rect 5707 10914 5735 10980
tri 5735 10914 5801 10980 sw
tri 6161 10972 6169 10980 ne
rect 6169 10972 6391 10980
tri 6169 10914 6227 10972 ne
rect 6227 10914 6391 10972
rect 4787 10907 5622 10914
rect 4368 10906 4701 10907
rect 0 10821 4283 10906
tri 4283 10821 4368 10906 sw
tri 4368 10821 4453 10906 ne
rect 4453 10821 4701 10906
tri 4701 10821 4787 10907 sw
tri 4787 10821 4873 10907 ne
rect 4873 10886 5622 10907
tri 5622 10886 5650 10914 sw
tri 5707 10886 5735 10914 ne
rect 5735 10886 5801 10914
tri 5801 10886 5829 10914 sw
tri 6227 10886 6255 10914 ne
rect 6255 10886 6391 10914
rect 4873 10821 5650 10886
rect 0 10813 4368 10821
tri 4368 10813 4376 10821 sw
tri 4453 10813 4461 10821 ne
rect 4461 10814 4787 10821
tri 4787 10814 4794 10821 sw
tri 4873 10814 4880 10821 ne
rect 4880 10814 5650 10821
rect 4461 10813 4794 10814
rect 0 10728 4376 10813
tri 4376 10728 4461 10813 sw
tri 4461 10728 4546 10813 ne
rect 4546 10728 4794 10813
tri 4794 10728 4880 10814 sw
tri 4880 10728 4966 10814 ne
rect 4966 10801 5650 10814
tri 5650 10801 5735 10886 sw
tri 5735 10801 5820 10886 ne
rect 5820 10801 5829 10886
rect 4966 10792 5735 10801
tri 5735 10792 5744 10801 sw
tri 5820 10792 5829 10801 ne
tri 5829 10792 5923 10886 sw
tri 6255 10885 6256 10886 ne
rect 6256 10885 6391 10886
rect 6627 11026 6800 11121
rect 7036 11028 7101 11262
tri 7101 11028 7375 11302 sw
tri 7489 11292 7499 11302 ne
rect 7499 11292 7598 11302
rect 7834 11428 8009 11528
rect 8245 11428 8250 11664
rect 7834 11415 8250 11428
tri 8250 11415 8637 11802 sw
tri 8637 11415 9024 11802 ne
rect 9024 11771 10191 11802
rect 10427 12004 12226 12007
rect 12462 12215 14683 12240
rect 12462 12191 13547 12215
rect 12462 12004 12923 12191
rect 10427 11976 12923 12004
rect 10427 11771 10870 11976
rect 9024 11740 10870 11771
rect 11106 11955 12923 11976
rect 13159 11979 13547 12191
rect 13783 12170 14683 12215
rect 13783 11979 14244 12170
rect 13159 11955 14244 11979
rect 11106 11934 14244 11955
rect 14480 12155 14683 12170
tri 14683 12155 15342 12814 sw
rect 35157 12734 35250 12970
rect 35486 12734 35584 12970
rect 35820 12734 35918 12970
rect 36154 12734 36252 12970
rect 36488 12734 36586 12970
rect 36822 12734 36920 12970
rect 37156 12734 37254 12970
rect 37490 12734 37588 12970
rect 37824 12734 37922 12970
rect 38158 12734 38256 12970
rect 38492 12734 38590 12970
rect 38826 12734 38924 12970
rect 39160 12734 39258 12970
rect 39494 12734 39592 12970
rect 39828 12734 40000 12970
rect 35157 12648 40000 12734
rect 35157 12412 35250 12648
rect 35486 12412 35584 12648
rect 35820 12412 35918 12648
rect 36154 12412 36252 12648
rect 36488 12412 36586 12648
rect 36822 12412 36920 12648
rect 37156 12412 37254 12648
rect 37490 12412 37588 12648
rect 37824 12412 37922 12648
rect 38158 12412 38256 12648
rect 38492 12412 38590 12648
rect 38826 12412 38924 12648
rect 39160 12412 39258 12648
rect 39494 12412 39592 12648
rect 39828 12412 40000 12648
rect 35157 12326 40000 12412
rect 14480 11934 14903 12155
rect 11106 11927 14903 11934
rect 11106 11740 11567 11927
rect 9024 11732 11567 11740
rect 9024 11496 9494 11732
rect 9730 11691 11567 11732
rect 11803 11919 14903 11927
rect 15139 11919 15342 12155
rect 11803 11916 15342 11919
rect 11803 11691 12226 11916
rect 9730 11683 12226 11691
rect 9730 11496 10191 11683
rect 9024 11447 10191 11496
rect 10427 11680 12226 11683
rect 12462 11891 15342 11916
rect 12462 11867 13547 11891
rect 12462 11680 12923 11867
rect 10427 11652 12923 11680
rect 10427 11447 10870 11652
rect 9024 11416 10870 11447
rect 11106 11631 12923 11652
rect 13159 11655 13547 11867
rect 13783 11848 15342 11891
rect 13783 11655 14244 11848
rect 13159 11631 14244 11655
rect 11106 11612 14244 11631
rect 14480 11834 15342 11848
rect 14480 11612 14903 11834
rect 11106 11603 14903 11612
rect 11106 11416 11567 11603
rect 9024 11415 11567 11416
rect 7834 11292 8637 11415
tri 7499 11028 7763 11292 ne
rect 7763 11260 8637 11292
tri 8637 11260 8792 11415 sw
tri 9024 11260 9179 11415 ne
rect 9179 11407 11567 11415
rect 9179 11260 9494 11407
rect 7763 11117 8413 11260
rect 7763 11028 8009 11117
rect 7036 11026 7375 11028
rect 6627 10914 7375 11026
tri 7375 10914 7489 11028 sw
tri 7763 10914 7877 11028 ne
rect 7877 10914 8009 11028
rect 6627 10898 7489 10914
rect 6627 10885 7161 10898
tri 6256 10792 6349 10885 ne
rect 6349 10792 7161 10885
rect 4966 10728 5744 10792
rect 0 10643 4461 10728
tri 4461 10643 4546 10728 sw
tri 4546 10643 4631 10728 ne
rect 4631 10643 4880 10728
rect 0 10568 4546 10643
tri 4546 10568 4621 10643 sw
tri 4631 10568 4706 10643 ne
rect 4706 10642 4880 10643
tri 4880 10642 4966 10728 sw
tri 4966 10642 5052 10728 ne
rect 5052 10707 5744 10728
tri 5744 10707 5829 10792 sw
tri 5829 10707 5914 10792 ne
rect 5914 10707 5923 10792
rect 5052 10698 5829 10707
tri 5829 10698 5838 10707 sw
tri 5914 10698 5923 10707 ne
tri 5923 10698 6017 10792 sw
tri 6349 10698 6443 10792 ne
rect 6443 10715 7161 10792
rect 6443 10698 6800 10715
rect 5052 10642 5838 10698
rect 4706 10569 4966 10642
tri 4966 10569 5039 10642 sw
tri 5052 10569 5125 10642 ne
rect 5125 10613 5838 10642
tri 5838 10613 5923 10698 sw
tri 5923 10613 6008 10698 ne
rect 6008 10613 6017 10698
rect 5125 10604 5923 10613
tri 5923 10604 5932 10613 sw
tri 6008 10604 6017 10613 ne
tri 6017 10604 6111 10698 sw
tri 6443 10604 6537 10698 ne
rect 6537 10604 6800 10698
rect 5125 10569 5932 10604
rect 4706 10568 5039 10569
rect 0 10483 4621 10568
tri 4621 10483 4706 10568 sw
tri 4706 10483 4791 10568 ne
rect 4791 10483 5039 10568
tri 5039 10483 5125 10569 sw
tri 5125 10483 5211 10569 ne
rect 5211 10519 5932 10569
tri 5932 10519 6017 10604 sw
tri 6017 10519 6102 10604 ne
rect 6102 10546 6111 10604
tri 6111 10546 6169 10604 sw
tri 6537 10546 6595 10604 ne
rect 6595 10546 6800 10604
rect 6102 10519 6169 10546
rect 5211 10510 6017 10519
tri 6017 10510 6026 10519 sw
tri 6102 10510 6111 10519 ne
rect 6111 10510 6169 10519
tri 6169 10510 6205 10546 sw
tri 6595 10510 6631 10546 ne
rect 6631 10510 6800 10546
rect 5211 10483 6026 10510
rect 0 10479 4706 10483
tri 4706 10479 4710 10483 sw
tri 4791 10479 4795 10483 ne
rect 4795 10480 5125 10483
tri 5125 10480 5128 10483 sw
tri 5211 10480 5214 10483 ne
rect 5214 10480 6026 10483
rect 4795 10479 5128 10480
rect 0 10406 4710 10479
tri 3940 10346 4000 10406 ne
rect 4000 10394 4710 10406
tri 4710 10394 4795 10479 sw
tri 4795 10394 4880 10479 ne
rect 4880 10394 5128 10479
tri 5128 10394 5214 10480 sw
tri 5214 10394 5300 10480 ne
rect 5300 10452 6026 10480
tri 6026 10452 6084 10510 sw
tri 6111 10452 6169 10510 ne
rect 6169 10452 6205 10510
rect 5300 10416 6084 10452
tri 6084 10416 6120 10452 sw
tri 6169 10416 6205 10452 ne
tri 6205 10416 6299 10510 sw
tri 6631 10416 6725 10510 ne
rect 6725 10479 6800 10510
rect 7036 10662 7161 10715
rect 7397 10662 7489 10898
rect 7036 10526 7489 10662
tri 7489 10526 7877 10914 sw
tri 7877 10881 7910 10914 ne
rect 7910 10881 8009 10914
rect 8245 11024 8413 11117
rect 8649 11028 8792 11260
tri 8792 11028 9024 11260 sw
tri 9179 11028 9411 11260 ne
rect 9411 11171 9494 11260
rect 9730 11367 11567 11407
rect 11803 11598 14903 11603
rect 15139 11598 15342 11834
rect 11803 11592 15342 11598
rect 11803 11367 12226 11592
rect 9730 11359 12226 11367
rect 9730 11171 10191 11359
rect 9411 11123 10191 11171
rect 10427 11356 12226 11359
rect 12462 11567 15342 11592
rect 12462 11543 13547 11567
rect 12462 11356 12923 11543
rect 10427 11328 12923 11356
rect 10427 11123 10870 11328
rect 9411 11092 10870 11123
rect 11106 11307 12923 11328
rect 13159 11331 13547 11543
rect 13783 11526 15342 11567
rect 13783 11331 14244 11526
rect 13159 11307 14244 11331
rect 11106 11290 14244 11307
rect 14480 11513 15342 11526
rect 14480 11290 14903 11513
rect 11106 11279 14903 11290
rect 11106 11092 11567 11279
rect 9411 11043 11567 11092
rect 11803 11277 14903 11279
rect 15139 11458 15342 11513
tri 15342 11458 16039 12155 sw
rect 35157 12090 35250 12326
rect 35486 12090 35584 12326
rect 35820 12090 35918 12326
rect 36154 12090 36252 12326
rect 36488 12090 36586 12326
rect 36822 12090 36920 12326
rect 37156 12090 37254 12326
rect 37490 12090 37588 12326
rect 37824 12090 37922 12326
rect 38158 12090 38256 12326
rect 38492 12090 38590 12326
rect 38826 12090 38924 12326
rect 39160 12090 39258 12326
rect 39494 12090 39592 12326
rect 39828 12090 40000 12326
rect 35157 12004 40000 12090
rect 35157 11768 35250 12004
rect 35486 11768 35584 12004
rect 35820 11768 35918 12004
rect 36154 11768 36252 12004
rect 36488 11768 36586 12004
rect 36822 11768 36920 12004
rect 37156 11768 37254 12004
rect 37490 11768 37588 12004
rect 37824 11768 37922 12004
rect 38158 11768 38256 12004
rect 38492 11768 38590 12004
rect 38826 11768 38924 12004
rect 39160 11768 39258 12004
rect 39494 11768 39592 12004
rect 39828 11768 40000 12004
rect 35157 11682 40000 11768
rect 15139 11277 15600 11458
rect 11803 11268 15600 11277
rect 11803 11043 12226 11268
rect 9411 11035 12226 11043
rect 9411 11028 10191 11035
rect 8649 11024 9024 11028
rect 8245 10881 9024 11024
tri 7910 10526 8265 10881 ne
rect 8265 10861 9024 10881
tri 9024 10861 9191 11028 sw
tri 9411 10861 9578 11028 ne
rect 9578 10861 10191 11028
rect 8265 10713 8812 10861
rect 8265 10526 8413 10713
rect 7036 10494 7877 10526
rect 7036 10479 7565 10494
rect 6725 10416 7565 10479
rect 5300 10394 6120 10416
rect 4000 10367 4795 10394
tri 4795 10367 4822 10394 sw
tri 4880 10367 4907 10394 ne
rect 4907 10367 5214 10394
tri 5214 10367 5241 10394 sw
tri 5300 10367 5327 10394 ne
rect 5327 10367 6120 10394
tri 6120 10367 6169 10416 sw
tri 6205 10367 6254 10416 ne
rect 6254 10367 6299 10416
tri 6299 10367 6348 10416 sw
tri 6725 10367 6774 10416 ne
rect 6774 10367 7565 10416
rect 4000 10346 4822 10367
rect 0 10280 3915 10346
tri 3915 10280 3981 10346 sw
tri 4000 10280 4066 10346 ne
rect 4066 10309 4822 10346
tri 4822 10309 4880 10367 sw
tri 4907 10309 4965 10367 ne
rect 4965 10309 5241 10367
rect 4066 10280 4880 10309
tri 3887 10186 3981 10280 ne
tri 3981 10271 3990 10280 sw
tri 4066 10271 4075 10280 ne
rect 4075 10271 4880 10280
rect 3981 10186 3990 10271
tri 3990 10186 4075 10271 sw
tri 4075 10186 4160 10271 ne
rect 4160 10224 4880 10271
tri 4880 10224 4965 10309 sw
tri 4965 10224 5050 10309 ne
rect 5050 10281 5241 10309
tri 5241 10281 5327 10367 sw
tri 5327 10281 5413 10367 ne
rect 5413 10322 6169 10367
tri 6169 10322 6214 10367 sw
tri 6254 10322 6299 10367 ne
rect 6299 10322 6348 10367
tri 6348 10322 6393 10367 sw
tri 6774 10322 6819 10367 ne
rect 6819 10351 7565 10367
rect 6819 10322 7161 10351
rect 5413 10281 6214 10322
rect 5050 10232 5327 10281
tri 5327 10232 5376 10281 sw
tri 5413 10232 5462 10281 ne
rect 5462 10237 6214 10281
tri 6214 10237 6299 10322 sw
tri 6299 10237 6384 10322 ne
rect 6384 10237 6393 10322
rect 5462 10232 6299 10237
rect 5050 10224 5376 10232
rect 4160 10186 4965 10224
tri 3981 10092 4075 10186 ne
tri 4075 10177 4084 10186 sw
tri 4160 10177 4169 10186 ne
rect 4169 10177 4965 10186
rect 4075 10092 4084 10177
tri 4084 10092 4169 10177 sw
tri 4169 10092 4254 10177 ne
rect 4254 10145 4965 10177
tri 4965 10145 5044 10224 sw
tri 5050 10145 5129 10224 ne
rect 5129 10146 5376 10224
tri 5376 10146 5462 10232 sw
tri 5462 10146 5548 10232 ne
rect 5548 10228 6299 10232
tri 6299 10228 6308 10237 sw
tri 6384 10228 6393 10237 ne
tri 6393 10228 6487 10322 sw
tri 6819 10228 6913 10322 ne
rect 6913 10228 7161 10322
rect 5548 10146 6308 10228
rect 5129 10145 5462 10146
rect 4254 10092 5044 10145
tri 4075 9998 4169 10092 ne
tri 4169 10083 4178 10092 sw
tri 4254 10083 4263 10092 ne
rect 4263 10083 5044 10092
rect 4169 9998 4178 10083
tri 4178 9998 4263 10083 sw
tri 4263 9998 4348 10083 ne
rect 4348 10060 5044 10083
tri 5044 10060 5129 10145 sw
tri 5129 10060 5214 10145 ne
rect 5214 10060 5462 10145
tri 5462 10060 5548 10146 sw
tri 5548 10060 5634 10146 ne
rect 5634 10143 6308 10146
tri 6308 10143 6393 10228 sw
tri 6393 10143 6478 10228 ne
rect 6478 10143 6487 10228
rect 5634 10134 6393 10143
tri 6393 10134 6402 10143 sw
tri 6478 10134 6487 10143 ne
tri 6487 10134 6581 10228 sw
tri 6913 10134 7007 10228 ne
rect 7007 10134 7161 10228
rect 5634 10060 6402 10134
rect 4348 9998 5129 10060
tri 4169 9980 4187 9998 ne
rect 4187 9989 4263 9998
tri 4263 9989 4272 9998 sw
tri 4348 9989 4357 9998 ne
rect 4357 9989 5129 9998
rect 4187 9980 4272 9989
tri 4272 9980 4281 9989 sw
tri 4357 9980 4366 9989 ne
rect 4366 9980 5129 9989
rect 0 9978 3764 9980
tri 3764 9978 3766 9980 sw
tri 4187 9978 4189 9980 ne
rect 4189 9978 4281 9980
tri 4281 9978 4283 9980 sw
tri 4366 9978 4368 9980 ne
rect 4368 9978 5129 9980
tri 5129 9978 5211 10060 sw
tri 5214 9978 5296 10060 ne
rect 5296 9978 5548 10060
tri 5548 9978 5630 10060 sw
tri 5634 9978 5716 10060 ne
rect 5716 10049 6402 10060
tri 6402 10049 6487 10134 sw
tri 6487 10049 6572 10134 ne
rect 6572 10049 6581 10134
rect 5716 10040 6487 10049
tri 6487 10040 6496 10049 sw
tri 6572 10040 6581 10049 ne
tri 6581 10040 6675 10134 sw
tri 7007 10130 7011 10134 ne
rect 7011 10130 7161 10134
tri 7011 10040 7101 10130 ne
rect 7101 10115 7161 10130
rect 7397 10258 7565 10351
rect 7801 10428 7877 10494
tri 7877 10428 7975 10526 sw
tri 8265 10428 8363 10526 ne
rect 8363 10477 8413 10526
rect 8649 10625 8812 10713
rect 9048 10641 9191 10861
tri 9191 10641 9411 10861 sw
tri 9578 10641 9798 10861 ne
rect 9798 10799 10191 10861
rect 10427 11032 12226 11035
rect 12462 11243 15600 11268
rect 12462 11219 13547 11243
rect 12462 11032 12923 11219
rect 10427 11004 12923 11032
rect 10427 10799 10870 11004
rect 9798 10768 10870 10799
rect 11106 10983 12923 11004
rect 13159 11007 13547 11219
rect 13783 11222 15600 11243
rect 15836 11222 16039 11458
rect 13783 11204 16039 11222
rect 13783 11007 14244 11204
rect 13159 10983 14244 11007
rect 11106 10968 14244 10983
rect 14480 11192 16039 11204
rect 14480 10968 14903 11192
rect 11106 10956 14903 10968
rect 15139 11127 16039 11192
rect 15139 10956 15600 11127
rect 11106 10955 15600 10956
rect 11106 10768 11567 10955
rect 9798 10719 11567 10768
rect 11803 10944 15600 10955
rect 11803 10719 12226 10944
rect 9798 10710 12226 10719
rect 9798 10641 10191 10710
rect 9048 10625 9411 10641
rect 8649 10541 9411 10625
tri 9411 10541 9511 10641 sw
tri 9798 10541 9898 10641 ne
rect 9898 10541 10191 10641
rect 8649 10477 9511 10541
rect 8363 10457 9511 10477
rect 8363 10428 9216 10457
rect 7801 10258 7975 10428
rect 7397 10115 7975 10258
rect 7101 10088 7975 10115
tri 7975 10088 8315 10428 sw
tri 8363 10088 8703 10428 ne
rect 8703 10314 9216 10428
rect 8703 10088 8812 10314
rect 7101 10040 7971 10088
rect 5716 9978 6496 10040
rect 0 9920 3766 9978
rect 0 9684 295 9920
rect 531 9684 830 9920
rect 1066 9684 1365 9920
rect 1601 9684 1900 9920
rect 2136 9684 2434 9920
rect 2670 9684 2968 9920
rect 3204 9684 3502 9920
rect 3738 9793 3766 9920
tri 3766 9793 3951 9978 sw
tri 4189 9904 4263 9978 ne
rect 4263 9904 4283 9978
tri 4283 9904 4357 9978 sw
tri 4368 9904 4442 9978 ne
rect 4442 9975 5211 9978
tri 5211 9975 5214 9978 sw
tri 5296 9975 5299 9978 ne
rect 5299 9975 5630 9978
rect 4442 9904 5214 9975
tri 4263 9810 4357 9904 ne
tri 4357 9895 4366 9904 sw
tri 4442 9895 4451 9904 ne
rect 4451 9895 5214 9904
rect 4357 9810 4366 9895
tri 4366 9810 4451 9895 sw
tri 4451 9810 4536 9895 ne
rect 4536 9890 5214 9895
tri 5214 9890 5299 9975 sw
tri 5299 9890 5384 9975 ne
rect 5384 9892 5630 9975
tri 5630 9892 5716 9978 sw
tri 5716 9892 5802 9978 ne
rect 5802 9955 6496 9978
tri 6496 9955 6581 10040 sw
tri 6581 9955 6666 10040 ne
rect 6666 9955 6675 10040
rect 5802 9946 6581 9955
tri 6581 9946 6590 9955 sw
tri 6666 9946 6675 9955 ne
tri 6675 9946 6769 10040 sw
tri 7101 9946 7195 10040 ne
rect 7195 9947 7971 10040
rect 7195 9946 7565 9947
rect 5802 9892 6590 9946
rect 5384 9890 5716 9892
rect 4536 9878 5299 9890
tri 5299 9878 5311 9890 sw
tri 5384 9878 5396 9890 ne
rect 5396 9878 5716 9890
rect 4536 9810 5311 9878
tri 4357 9793 4374 9810 ne
rect 4374 9801 4451 9810
tri 4451 9801 4460 9810 sw
tri 4536 9801 4545 9810 ne
rect 4545 9801 5311 9810
rect 4374 9793 4460 9801
tri 4460 9793 4468 9801 sw
tri 4545 9793 4553 9801 ne
rect 4553 9793 5311 9801
tri 5311 9793 5396 9878 sw
tri 5396 9793 5481 9878 ne
rect 5481 9812 5716 9878
tri 5716 9812 5796 9892 sw
tri 5802 9812 5882 9892 ne
rect 5882 9861 6590 9892
tri 6590 9861 6675 9946 sw
tri 6675 9861 6760 9946 ne
rect 6760 9861 6769 9946
rect 5882 9852 6675 9861
tri 6675 9852 6684 9861 sw
tri 6760 9852 6769 9861 ne
tri 6769 9852 6863 9946 sw
tri 7195 9852 7289 9946 ne
rect 7289 9852 7565 9946
rect 5882 9812 6684 9852
rect 5481 9793 5796 9812
rect 3738 9716 3951 9793
tri 3951 9716 4028 9793 sw
tri 4374 9716 4451 9793 ne
rect 4451 9716 4468 9793
tri 4468 9716 4545 9793 sw
tri 4553 9716 4630 9793 ne
rect 4630 9726 5396 9793
tri 5396 9726 5463 9793 sw
tri 5481 9726 5548 9793 ne
rect 5548 9726 5796 9793
tri 5796 9726 5882 9812 sw
tri 5882 9726 5968 9812 ne
rect 5968 9767 6684 9812
tri 6684 9767 6769 9852 sw
tri 6769 9767 6854 9852 ne
rect 6854 9767 6863 9852
rect 5968 9758 6769 9767
tri 6769 9758 6778 9767 sw
tri 6854 9758 6863 9767 ne
tri 6863 9758 6957 9852 sw
tri 7289 9758 7383 9852 ne
rect 7383 9758 7565 9852
rect 5968 9726 6778 9758
rect 4630 9716 5463 9726
rect 3738 9684 4028 9716
rect 0 9622 4028 9684
tri 4028 9622 4122 9716 sw
tri 4451 9622 4545 9716 ne
tri 4545 9707 4554 9716 sw
tri 4630 9707 4639 9716 ne
rect 4639 9707 5463 9716
rect 4545 9622 4554 9707
tri 4554 9622 4639 9707 sw
tri 4639 9622 4724 9707 ne
rect 4724 9641 5463 9707
tri 5463 9641 5548 9726 sw
tri 5548 9641 5633 9726 ne
rect 5633 9641 5882 9726
rect 4724 9640 5548 9641
tri 5548 9640 5549 9641 sw
tri 5633 9640 5634 9641 ne
rect 5634 9640 5882 9641
tri 5882 9640 5968 9726 sw
tri 5968 9640 6054 9726 ne
rect 6054 9673 6778 9726
tri 6778 9673 6863 9758 sw
tri 6863 9673 6948 9758 ne
rect 6948 9704 6957 9758
tri 6957 9704 7011 9758 sw
tri 7383 9704 7437 9758 ne
rect 7437 9711 7565 9758
rect 7801 9852 7971 9947
rect 8207 10040 8315 10088
tri 8315 10040 8363 10088 sw
tri 8703 10040 8751 10088 ne
rect 8751 10078 8812 10088
rect 9048 10221 9216 10314
rect 9452 10221 9511 10457
rect 9048 10154 9511 10221
tri 9511 10154 9898 10541 sw
tri 9898 10474 9965 10541 ne
rect 9965 10474 10191 10541
rect 10427 10708 12226 10710
rect 12462 10919 15600 10944
rect 12462 10895 13547 10919
rect 12462 10708 12923 10895
rect 10427 10680 12923 10708
rect 10427 10474 10870 10680
tri 9965 10154 10285 10474 ne
rect 10285 10444 10870 10474
rect 11106 10659 12923 10680
rect 13159 10683 13547 10895
rect 13783 10891 15600 10919
rect 15836 11097 16039 11127
tri 16039 11097 16400 11458 sw
rect 35157 11446 35250 11682
rect 35486 11446 35584 11682
rect 35820 11446 35918 11682
rect 36154 11446 36252 11682
rect 36488 11446 36586 11682
rect 36822 11446 36920 11682
rect 37156 11446 37254 11682
rect 37490 11446 37588 11682
rect 37824 11446 37922 11682
rect 38158 11446 38256 11682
rect 38492 11446 38590 11682
rect 38826 11446 38924 11682
rect 39160 11446 39258 11682
rect 39494 11446 39592 11682
rect 39828 11446 40000 11682
rect 35157 11360 40000 11446
rect 35157 11124 35250 11360
rect 35486 11124 35584 11360
rect 35820 11124 35918 11360
rect 36154 11124 36252 11360
rect 36488 11124 36586 11360
rect 36822 11124 36920 11360
rect 37156 11124 37254 11360
rect 37490 11124 37588 11360
rect 37824 11124 37922 11360
rect 38158 11124 38256 11360
rect 38492 11124 38590 11360
rect 38826 11124 38924 11360
rect 39160 11124 39258 11360
rect 39494 11124 39592 11360
rect 39828 11124 40000 11360
rect 15836 10891 16073 11097
rect 13783 10882 16073 10891
rect 13783 10683 14244 10882
rect 13159 10659 14244 10683
rect 11106 10646 14244 10659
rect 14480 10871 16073 10882
rect 14480 10646 14903 10871
rect 11106 10635 14903 10646
rect 15139 10861 16073 10871
rect 16309 10861 16400 11097
rect 15139 10796 16400 10861
rect 15139 10635 15600 10796
rect 11106 10631 15600 10635
rect 11106 10444 11567 10631
rect 10285 10395 11567 10444
rect 11803 10620 15600 10631
rect 11803 10395 12226 10620
rect 10285 10384 12226 10395
rect 12462 10595 15600 10620
rect 12462 10571 13547 10595
rect 12462 10384 12923 10571
rect 10285 10356 12923 10384
rect 10285 10154 10870 10356
rect 9048 10078 9898 10154
rect 8751 10040 9898 10078
rect 8207 9852 8363 10040
rect 7801 9767 8363 9852
tri 8363 9767 8636 10040 sw
tri 8751 9767 9024 10040 ne
rect 9024 10024 9898 10040
rect 9024 9910 9649 10024
rect 9024 9767 9216 9910
rect 7801 9711 8636 9767
rect 7437 9704 8636 9711
rect 6948 9673 7011 9704
rect 6054 9664 6863 9673
tri 6863 9664 6872 9673 sw
tri 6948 9664 6957 9673 ne
rect 6957 9664 7011 9673
tri 7011 9664 7051 9704 sw
tri 7437 9664 7477 9704 ne
rect 7477 9697 8636 9704
rect 7477 9664 8365 9697
rect 6054 9652 6872 9664
tri 6872 9652 6884 9664 sw
tri 6957 9652 6969 9664 ne
rect 6969 9652 7051 9664
tri 7051 9652 7063 9664 sw
tri 7477 9652 7489 9664 ne
rect 7489 9652 8365 9664
rect 6054 9640 6884 9652
rect 4724 9622 5549 9640
rect 0 9541 4122 9622
rect 0 9346 3820 9541
rect 0 9110 295 9346
rect 531 9110 830 9346
rect 1066 9110 1365 9346
rect 1601 9110 1900 9346
rect 2136 9110 2434 9346
rect 2670 9110 2968 9346
rect 3204 9110 3502 9346
rect 3738 9305 3820 9346
rect 4056 9528 4122 9541
tri 4122 9528 4216 9622 sw
tri 4545 9528 4639 9622 ne
tri 4639 9613 4648 9622 sw
tri 4724 9613 4733 9622 ne
rect 4733 9613 5549 9622
rect 4639 9528 4648 9613
tri 4648 9528 4733 9613 sw
tri 4733 9528 4818 9613 ne
rect 4818 9610 5549 9613
tri 5549 9610 5579 9640 sw
tri 5634 9610 5664 9640 ne
rect 5664 9610 5968 9640
rect 4818 9528 5579 9610
rect 4056 9305 4216 9528
rect 3738 9191 4216 9305
tri 4216 9191 4553 9528 sw
tri 4639 9434 4733 9528 ne
tri 4733 9519 4742 9528 sw
tri 4818 9519 4827 9528 ne
rect 4827 9525 5579 9528
tri 5579 9525 5664 9610 sw
tri 5664 9525 5749 9610 ne
rect 5749 9554 5968 9610
tri 5968 9554 6054 9640 sw
tri 6054 9554 6140 9640 ne
rect 6140 9610 6884 9640
tri 6884 9610 6926 9652 sw
tri 6969 9610 7011 9652 ne
rect 7011 9610 7063 9652
rect 6140 9570 6926 9610
tri 6926 9570 6966 9610 sw
tri 7011 9570 7051 9610 ne
rect 7051 9570 7063 9610
tri 7063 9570 7145 9652 sw
tri 7489 9570 7571 9652 ne
rect 7571 9570 8365 9652
rect 6140 9554 6966 9570
rect 5749 9525 6054 9554
tri 6054 9525 6083 9554 sw
tri 6140 9525 6169 9554 ne
rect 6169 9525 6966 9554
tri 6966 9525 7011 9570 sw
tri 7051 9525 7096 9570 ne
rect 7096 9525 7145 9570
tri 7145 9525 7190 9570 sw
tri 7571 9525 7616 9570 ne
rect 7616 9541 8365 9570
rect 7616 9525 7971 9541
rect 4827 9519 5664 9525
rect 4733 9434 4742 9519
tri 4742 9434 4827 9519 sw
tri 4827 9434 4912 9519 ne
rect 4912 9477 5664 9519
tri 5664 9477 5712 9525 sw
tri 5749 9477 5797 9525 ne
rect 5797 9478 6083 9525
tri 6083 9478 6130 9525 sw
tri 6169 9478 6216 9525 ne
rect 6216 9478 7011 9525
rect 5797 9477 6130 9478
rect 4912 9434 5712 9477
tri 4733 9340 4827 9434 ne
tri 4827 9425 4836 9434 sw
tri 4912 9425 4921 9434 ne
rect 4921 9425 5712 9434
rect 4827 9340 4836 9425
tri 4836 9340 4921 9425 sw
tri 4921 9340 5006 9425 ne
rect 5006 9392 5712 9425
tri 5712 9392 5797 9477 sw
tri 5797 9392 5882 9477 ne
rect 5882 9392 6130 9477
tri 6130 9392 6216 9478 sw
tri 6216 9392 6302 9478 ne
rect 6302 9476 7011 9478
tri 7011 9476 7060 9525 sw
tri 7096 9476 7145 9525 ne
rect 7145 9476 7190 9525
tri 7190 9476 7239 9525 sw
tri 7616 9476 7665 9525 ne
rect 7665 9476 7971 9525
rect 6302 9392 7060 9476
rect 5006 9340 5797 9392
tri 4827 9246 4921 9340 ne
tri 4921 9331 4930 9340 sw
tri 5006 9331 5015 9340 ne
rect 5015 9331 5797 9340
rect 4921 9246 4930 9331
tri 4930 9246 5015 9331 sw
tri 5015 9246 5100 9331 ne
rect 5100 9307 5797 9331
tri 5797 9307 5882 9392 sw
tri 5882 9307 5967 9392 ne
rect 5967 9307 6216 9392
rect 5100 9246 5882 9307
tri 4921 9191 4976 9246 ne
rect 4976 9237 5015 9246
tri 5015 9237 5024 9246 sw
tri 5100 9237 5109 9246 ne
rect 5109 9237 5882 9246
rect 4976 9191 5024 9237
tri 5024 9191 5070 9237 sw
tri 5109 9191 5155 9237 ne
rect 5155 9222 5882 9237
tri 5882 9222 5967 9307 sw
tri 5967 9222 6052 9307 ne
rect 6052 9306 6216 9307
tri 6216 9306 6302 9392 sw
tri 6302 9306 6388 9392 ne
rect 6388 9391 7060 9392
tri 7060 9391 7145 9476 sw
tri 7145 9391 7230 9476 ne
rect 7230 9391 7239 9476
rect 6388 9382 7145 9391
tri 7145 9382 7154 9391 sw
tri 7230 9382 7239 9391 ne
tri 7239 9382 7333 9476 sw
tri 7665 9382 7759 9476 ne
rect 7759 9382 7971 9476
rect 6388 9306 7154 9382
rect 6052 9230 6302 9306
tri 6302 9230 6378 9306 sw
tri 6388 9230 6464 9306 ne
rect 6464 9297 7154 9306
tri 7154 9297 7239 9382 sw
tri 7239 9297 7324 9382 ne
rect 7324 9297 7333 9382
rect 6464 9288 7239 9297
tri 7239 9288 7248 9297 sw
tri 7324 9288 7333 9297 ne
tri 7333 9288 7427 9382 sw
tri 7759 9288 7853 9382 ne
rect 7853 9305 7971 9382
rect 8207 9461 8365 9541
rect 8601 9652 8636 9697
tri 8636 9652 8751 9767 sw
tri 9024 9652 9139 9767 ne
rect 9139 9674 9216 9767
rect 9452 9788 9649 9910
rect 9885 9788 9898 10024
rect 9452 9767 9898 9788
tri 9898 9767 10285 10154 sw
tri 10285 9767 10672 10154 ne
rect 10672 10120 10870 10154
rect 11106 10335 12923 10356
rect 13159 10359 13547 10571
rect 13783 10560 15600 10595
rect 15836 10560 16400 10796
rect 13783 10359 14244 10560
rect 13159 10335 14244 10359
rect 11106 10324 14244 10335
rect 14480 10550 16400 10560
rect 14480 10324 14903 10550
rect 11106 10314 14903 10324
rect 15139 10465 16400 10550
rect 15139 10314 15600 10465
rect 11106 10307 15600 10314
rect 11106 10120 11567 10307
rect 10672 10071 11567 10120
rect 11803 10296 15600 10307
rect 11803 10071 12226 10296
rect 10672 10060 12226 10071
rect 12462 10271 15600 10296
rect 12462 10247 13547 10271
rect 12462 10060 12923 10247
rect 10672 10031 12923 10060
rect 10672 9795 10870 10031
rect 11106 10011 12923 10031
rect 13159 10035 13547 10247
rect 13783 10238 15600 10271
rect 13783 10035 14244 10238
rect 13159 10011 14244 10035
rect 11106 10002 14244 10011
rect 14480 10229 15600 10238
rect 15836 10462 16400 10465
rect 15836 10229 16073 10462
rect 14480 10002 14903 10229
rect 11106 9993 14903 10002
rect 15139 10226 16073 10229
rect 16309 10226 16400 10462
rect 15139 10168 16400 10226
tri 16400 10168 17329 11097 sw
rect 35157 11038 40000 11124
rect 35157 10802 35250 11038
rect 35486 10802 35584 11038
rect 35820 10802 35918 11038
rect 36154 10802 36252 11038
rect 36488 10802 36586 11038
rect 36822 10802 36920 11038
rect 37156 10802 37254 11038
rect 37490 10802 37588 11038
rect 37824 10802 37922 11038
rect 38158 10802 38256 11038
rect 38492 10802 38590 11038
rect 38826 10802 38924 11038
rect 39160 10802 39258 11038
rect 39494 10802 39592 11038
rect 39828 10802 40000 11038
rect 35157 10716 40000 10802
rect 35157 10480 35250 10716
rect 35486 10480 35584 10716
rect 35820 10480 35918 10716
rect 36154 10480 36252 10716
rect 36488 10480 36586 10716
rect 36822 10480 36920 10716
rect 37156 10480 37254 10716
rect 37490 10480 37588 10716
rect 37824 10480 37922 10716
rect 38158 10480 38256 10716
rect 38492 10480 38590 10716
rect 38826 10480 38924 10716
rect 39160 10480 39258 10716
rect 39494 10480 39592 10716
rect 39828 10480 40000 10716
rect 35157 10394 40000 10480
rect 15139 10134 17329 10168
rect 15139 9993 15600 10134
rect 11106 9983 15600 9993
rect 11106 9795 11567 9983
rect 10672 9767 11567 9795
rect 9452 9674 10285 9767
rect 9139 9652 10285 9674
rect 8601 9461 8751 9652
rect 8207 9333 8751 9461
tri 8751 9333 9070 9652 sw
tri 9139 9333 9458 9652 ne
rect 9458 9620 10285 9652
tri 10285 9620 10432 9767 sw
tri 10672 9620 10819 9767 ne
rect 10819 9747 11567 9767
rect 11803 9972 15600 9983
rect 11803 9747 12226 9972
rect 10819 9736 12226 9747
rect 12462 9947 15600 9972
rect 12462 9923 13547 9947
rect 12462 9736 12923 9923
rect 10819 9687 12923 9736
rect 13159 9711 13547 9923
rect 13783 9915 15600 9947
rect 13783 9711 14244 9915
rect 13159 9687 14244 9711
rect 10819 9679 14244 9687
rect 14480 9908 15600 9915
rect 14480 9679 14903 9908
rect 10819 9672 14903 9679
rect 15139 9898 15600 9908
rect 15836 10079 17329 10134
rect 15836 9898 16050 10079
rect 15139 9843 16050 9898
rect 16286 9843 16545 10079
rect 16781 9843 17039 10079
rect 17275 9843 17329 10079
rect 15139 9803 17329 9843
rect 15139 9672 15600 9803
rect 10819 9659 15600 9672
rect 10819 9620 11567 9659
rect 9458 9477 10053 9620
rect 9458 9333 9649 9477
rect 8207 9305 8726 9333
rect 7853 9288 8726 9305
rect 6464 9230 7248 9288
rect 6052 9222 6378 9230
rect 5155 9220 5967 9222
tri 5967 9220 5969 9222 sw
tri 6052 9220 6054 9222 ne
rect 6054 9220 6378 9222
rect 5155 9191 5969 9220
rect 3738 9182 4553 9191
rect 3738 9110 4195 9182
rect 0 9050 4195 9110
tri 3370 8770 3650 9050 ne
rect 3650 8994 4195 9050
rect 3650 8770 3820 8994
rect 0 8702 3268 8770
rect 0 8466 267 8702
rect 503 8466 816 8702
rect 1052 8466 1365 8702
rect 1601 8466 1914 8702
rect 2150 8466 2463 8702
rect 2699 8466 3012 8702
rect 3248 8668 3268 8702
tri 3268 8668 3370 8770 sw
tri 3650 8668 3752 8770 ne
rect 3752 8758 3820 8770
rect 4056 8946 4195 8994
rect 4431 9135 4553 9182
tri 4553 9135 4609 9191 sw
tri 4976 9152 5015 9191 ne
rect 5015 9152 5070 9191
tri 5070 9152 5109 9191 sw
tri 5155 9152 5194 9191 ne
rect 5194 9152 5969 9191
tri 5015 9135 5032 9152 ne
rect 5032 9143 5109 9152
tri 5109 9143 5118 9152 sw
tri 5194 9143 5203 9152 ne
rect 5203 9143 5969 9152
rect 5032 9135 5118 9143
tri 5118 9135 5126 9143 sw
tri 5203 9135 5211 9143 ne
rect 5211 9135 5969 9143
tri 5969 9135 6054 9220 sw
tri 6054 9135 6139 9220 ne
rect 6139 9144 6378 9220
tri 6378 9144 6464 9230 sw
tri 6464 9144 6550 9230 ne
rect 6550 9203 7248 9230
tri 7248 9203 7333 9288 sw
tri 7333 9203 7418 9288 ne
rect 7418 9203 7427 9288
rect 6550 9194 7333 9203
tri 7333 9194 7342 9203 sw
tri 7418 9194 7427 9203 ne
tri 7427 9194 7521 9288 sw
tri 7853 9194 7947 9288 ne
rect 7947 9194 8726 9288
rect 6550 9144 7342 9194
rect 6139 9135 6464 9144
tri 6464 9135 6473 9144 sw
tri 6550 9135 6559 9144 ne
rect 6559 9135 7342 9144
rect 4431 9071 4609 9135
tri 4609 9071 4673 9135 sw
tri 5032 9071 5096 9135 ne
rect 5096 9071 5126 9135
tri 5126 9071 5190 9135 sw
tri 5211 9071 5275 9135 ne
rect 5275 9071 6054 9135
rect 4431 8946 4673 9071
rect 4056 8818 4673 8946
tri 4673 8818 4926 9071 sw
tri 5096 9058 5109 9071 ne
rect 5109 9058 5190 9071
tri 5190 9058 5203 9071 sw
tri 5275 9058 5288 9071 ne
rect 5288 9058 6054 9071
tri 6054 9058 6131 9135 sw
tri 6139 9058 6216 9135 ne
rect 6216 9058 6473 9135
tri 6473 9058 6550 9135 sw
tri 6559 9058 6636 9135 ne
rect 6636 9109 7342 9135
tri 7342 9109 7427 9194 sw
tri 7427 9109 7512 9194 ne
rect 7512 9109 7521 9194
rect 6636 9100 7427 9109
tri 7427 9100 7436 9109 sw
tri 7512 9100 7521 9109 ne
tri 7521 9100 7615 9194 sw
tri 7947 9100 8041 9194 ne
rect 8041 9150 8726 9194
rect 8041 9100 8365 9150
rect 6636 9058 7436 9100
tri 5109 8964 5203 9058 ne
tri 5203 9049 5212 9058 sw
tri 5288 9049 5297 9058 ne
rect 5297 9049 6131 9058
rect 5203 8964 5212 9049
tri 5212 8964 5297 9049 sw
tri 5297 8964 5382 9049 ne
rect 5382 8973 6131 9049
tri 6131 8973 6216 9058 sw
tri 6216 8973 6301 9058 ne
rect 6301 8973 6550 9058
rect 5382 8964 6216 8973
tri 5203 8870 5297 8964 ne
tri 5297 8955 5306 8964 sw
tri 5382 8955 5391 8964 ne
rect 5391 8955 6216 8964
rect 5297 8870 5306 8955
tri 5306 8870 5391 8955 sw
tri 5391 8870 5476 8955 ne
rect 5476 8888 6216 8955
tri 6216 8888 6301 8973 sw
tri 6301 8888 6386 8973 ne
rect 6386 8972 6550 8973
tri 6550 8972 6636 9058 sw
tri 6636 8972 6722 9058 ne
rect 6722 9015 7436 9058
tri 7436 9015 7521 9100 sw
tri 7521 9015 7606 9100 ne
rect 7606 9015 7615 9100
rect 6722 9006 7521 9015
tri 7521 9006 7530 9015 sw
tri 7606 9006 7615 9015 ne
tri 7615 9006 7709 9100 sw
tri 8041 9006 8135 9100 ne
rect 8135 9006 8365 9100
rect 6722 8972 7530 9006
rect 6386 8896 6636 8972
tri 6636 8896 6712 8972 sw
tri 6722 8896 6798 8972 ne
rect 6798 8921 7530 8972
tri 7530 8921 7615 9006 sw
tri 7615 8921 7700 9006 ne
rect 7700 8921 7709 9006
rect 6798 8912 7615 8921
tri 7615 8912 7624 8921 sw
tri 7700 8912 7709 8921 ne
tri 7709 8912 7803 9006 sw
tri 8135 8912 8229 9006 ne
rect 8229 8914 8365 9006
rect 8601 9097 8726 9150
rect 8962 9264 9070 9333
tri 9070 9264 9139 9333 sw
tri 9458 9264 9527 9333 ne
rect 9527 9264 9649 9333
rect 8962 9166 9139 9264
tri 9139 9166 9237 9264 sw
tri 9527 9166 9625 9264 ne
rect 9625 9241 9649 9264
rect 9885 9384 10053 9477
rect 10289 9384 10432 9620
rect 9885 9380 10432 9384
tri 10432 9380 10672 9620 sw
tri 10819 9380 11059 9620 ne
rect 11059 9423 11567 9620
rect 11803 9648 15600 9659
rect 11803 9423 12226 9648
rect 11059 9412 12226 9423
rect 12462 9623 15600 9648
rect 12462 9599 13547 9623
rect 12462 9412 12923 9599
rect 11059 9380 12923 9412
rect 9885 9280 10672 9380
tri 10672 9280 10772 9380 sw
tri 11059 9280 11159 9380 ne
rect 11159 9363 12923 9380
rect 13159 9387 13547 9599
rect 13783 9592 15600 9623
rect 13783 9387 14244 9592
rect 13159 9363 14244 9387
rect 11159 9356 14244 9363
rect 14480 9587 15600 9592
rect 14480 9356 14903 9587
rect 11159 9351 14903 9356
rect 15139 9567 15600 9587
rect 15836 9600 17329 9803
tri 17329 9600 17897 10168 sw
rect 35157 10158 35250 10394
rect 35486 10158 35584 10394
rect 35820 10158 35918 10394
rect 36154 10158 36252 10394
rect 36488 10158 36586 10394
rect 36822 10158 36920 10394
rect 37156 10158 37254 10394
rect 37490 10158 37588 10394
rect 37824 10158 37922 10394
rect 38158 10158 38256 10394
rect 38492 10158 38590 10394
rect 38826 10158 38924 10394
rect 39160 10158 39258 10394
rect 39494 10158 39592 10394
rect 39828 10158 40000 10394
rect 35157 10072 40000 10158
rect 35157 9836 35250 10072
rect 35486 9836 35584 10072
rect 35820 9836 35918 10072
rect 36154 9836 36252 10072
rect 36488 9836 36586 10072
rect 36822 9836 36920 10072
rect 37156 9836 37254 10072
rect 37490 9836 37588 10072
rect 37824 9836 37922 10072
rect 38158 9836 38256 10072
rect 38492 9836 38590 10072
rect 38826 9836 38924 10072
rect 39160 9836 39258 10072
rect 39494 9836 39592 10072
rect 39828 9836 40000 10072
rect 35157 9750 40000 9836
rect 15836 9599 17897 9600
rect 15836 9567 16065 9599
rect 15139 9471 16065 9567
rect 15139 9351 15600 9471
rect 11159 9334 15600 9351
rect 11159 9280 11567 9334
rect 9885 9241 10772 9280
rect 9625 9221 10772 9241
rect 9625 9166 10452 9221
rect 8962 9097 9237 9166
rect 8601 8929 9237 9097
tri 9237 8929 9474 9166 sw
tri 9625 8929 9862 9166 ne
rect 9862 9073 10452 9166
rect 9862 8929 10053 9073
rect 8601 8914 9130 8929
rect 8229 8912 9130 8914
rect 6798 8896 7624 8912
rect 6386 8888 6712 8896
rect 5476 8882 6301 8888
tri 6301 8882 6307 8888 sw
tri 6386 8882 6392 8888 ne
rect 6392 8882 6712 8888
rect 5476 8870 6307 8882
tri 5297 8818 5349 8870 ne
rect 5349 8861 5391 8870
tri 5391 8861 5400 8870 sw
tri 5476 8861 5485 8870 ne
rect 5485 8861 6307 8870
rect 5349 8818 5400 8861
rect 4056 8758 4556 8818
rect 3752 8668 4556 8758
rect 3248 8469 3370 8668
tri 3370 8469 3569 8668 sw
tri 3752 8469 3951 8668 ne
rect 3951 8635 4556 8668
rect 3951 8469 4195 8635
rect 3248 8466 3569 8469
rect 0 8362 3569 8466
rect 0 8126 267 8362
rect 503 8126 816 8362
rect 1052 8126 1365 8362
rect 1601 8126 1914 8362
rect 2150 8126 2463 8362
rect 2699 8126 3012 8362
rect 3248 8292 3569 8362
tri 3569 8292 3746 8469 sw
tri 3951 8292 4128 8469 ne
rect 4128 8399 4195 8469
rect 4431 8582 4556 8635
rect 4792 8770 4926 8818
tri 4926 8770 4974 8818 sw
tri 5349 8776 5391 8818 ne
rect 5391 8776 5400 8818
tri 5400 8776 5485 8861 sw
tri 5485 8776 5570 8861 ne
rect 5570 8797 6307 8861
tri 6307 8797 6392 8882 sw
tri 6392 8797 6477 8882 ne
rect 6477 8810 6712 8882
tri 6712 8810 6798 8896 sw
tri 6798 8810 6884 8896 ne
rect 6884 8827 7624 8896
tri 7624 8827 7709 8912 sw
tri 7709 8827 7794 8912 ne
rect 7794 8862 7803 8912
tri 7803 8862 7853 8912 sw
tri 8229 8862 8279 8912 ne
rect 8279 8862 9130 8912
rect 7794 8827 7853 8862
rect 6884 8818 7709 8827
tri 7709 8818 7718 8827 sw
tri 7794 8818 7803 8827 ne
rect 7803 8818 7853 8827
tri 7853 8818 7897 8862 sw
tri 8279 8818 8323 8862 ne
rect 8323 8818 9130 8862
rect 6884 8810 7718 8818
rect 6477 8797 6798 8810
tri 6798 8797 6811 8810 sw
tri 6884 8797 6897 8810 ne
rect 6897 8797 7718 8810
rect 5570 8776 6392 8797
tri 5391 8770 5397 8776 ne
rect 5397 8770 5485 8776
rect 4792 8582 4974 8770
rect 4431 8469 4974 8582
tri 4974 8469 5275 8770 sw
tri 5397 8682 5485 8770 ne
tri 5485 8767 5494 8776 sw
tri 5570 8767 5579 8776 ne
rect 5579 8767 6392 8776
rect 5485 8682 5494 8767
tri 5494 8682 5579 8767 sw
tri 5579 8682 5664 8767 ne
rect 5664 8724 6392 8767
tri 6392 8724 6465 8797 sw
tri 6477 8724 6550 8797 ne
rect 6550 8724 6811 8797
tri 6811 8724 6884 8797 sw
tri 6897 8724 6970 8797 ne
rect 6970 8768 7718 8797
tri 7718 8768 7768 8818 sw
tri 7803 8768 7853 8818 ne
rect 7853 8768 7897 8818
rect 6970 8724 7768 8768
tri 7768 8724 7812 8768 sw
tri 7853 8724 7897 8768 ne
tri 7897 8724 7991 8818 sw
tri 8323 8724 8417 8818 ne
rect 8417 8786 9130 8818
rect 8417 8724 8726 8786
rect 5664 8683 6465 8724
tri 6465 8683 6506 8724 sw
tri 6550 8683 6591 8724 ne
rect 6591 8683 6884 8724
tri 6884 8683 6925 8724 sw
tri 6970 8683 7011 8724 ne
rect 7011 8683 7812 8724
tri 7812 8683 7853 8724 sw
tri 7897 8683 7938 8724 ne
rect 7938 8683 7991 8724
tri 7991 8683 8032 8724 sw
tri 8417 8683 8458 8724 ne
rect 8458 8683 8726 8724
rect 5664 8682 6506 8683
tri 5485 8588 5579 8682 ne
tri 5579 8673 5588 8682 sw
tri 5664 8673 5673 8682 ne
rect 5673 8673 6506 8682
rect 5579 8588 5588 8673
tri 5588 8588 5673 8673 sw
tri 5673 8588 5758 8673 ne
rect 5758 8639 6506 8673
tri 6506 8639 6550 8683 sw
tri 6591 8639 6635 8683 ne
rect 6635 8639 6925 8683
rect 5758 8588 6550 8639
tri 5579 8494 5673 8588 ne
tri 5673 8579 5682 8588 sw
tri 5758 8579 5767 8588 ne
rect 5767 8579 6550 8588
rect 5673 8494 5682 8579
tri 5682 8494 5767 8579 sw
tri 5767 8494 5852 8579 ne
rect 5852 8554 6550 8579
tri 6550 8554 6635 8639 sw
tri 6635 8554 6720 8639 ne
rect 6720 8597 6925 8639
tri 6925 8597 7011 8683 sw
tri 7011 8597 7097 8683 ne
rect 7097 8630 7853 8683
tri 7853 8630 7906 8683 sw
tri 7938 8630 7991 8683 ne
rect 7991 8630 8032 8683
tri 8032 8630 8085 8683 sw
tri 8458 8630 8511 8683 ne
rect 8511 8630 8726 8683
rect 7097 8597 7906 8630
rect 6720 8562 7011 8597
tri 7011 8562 7046 8597 sw
tri 7097 8562 7132 8597 ne
rect 7132 8562 7906 8597
rect 6720 8554 7046 8562
rect 5852 8494 6635 8554
tri 5673 8469 5698 8494 ne
rect 5698 8485 5767 8494
tri 5767 8485 5776 8494 sw
tri 5852 8485 5861 8494 ne
rect 5861 8485 6635 8494
rect 5698 8469 5776 8485
tri 5776 8469 5792 8485 sw
tri 5861 8469 5877 8485 ne
rect 5877 8469 6635 8485
tri 6635 8469 6720 8554 sw
tri 6720 8469 6805 8554 ne
rect 6805 8476 7046 8554
tri 7046 8476 7132 8562 sw
tri 7132 8476 7218 8562 ne
rect 7218 8545 7906 8562
tri 7906 8545 7991 8630 sw
tri 7991 8545 8076 8630 ne
rect 8076 8545 8085 8630
rect 7218 8536 7991 8545
tri 7991 8536 8000 8545 sw
tri 8076 8536 8085 8545 ne
tri 8085 8536 8179 8630 sw
tri 8511 8536 8605 8630 ne
rect 8605 8550 8726 8630
rect 8962 8693 9130 8786
rect 9366 8778 9474 8929
tri 9474 8778 9625 8929 sw
tri 9862 8778 10013 8929 ne
rect 10013 8837 10053 8929
rect 10289 8985 10452 9073
rect 10688 8985 10772 9221
rect 10289 8893 10772 8985
tri 10772 8893 11159 9280 sw
tri 11159 9098 11341 9280 ne
rect 11341 9098 11567 9280
rect 11803 9324 15600 9334
rect 11803 9098 12226 9324
tri 11341 8893 11546 9098 ne
rect 11546 9088 12226 9098
rect 12462 9299 15600 9324
rect 12462 9275 13547 9299
rect 12462 9088 12923 9275
rect 11546 9039 12923 9088
rect 13159 9063 13547 9275
rect 13783 9269 15600 9299
rect 13783 9063 14244 9269
rect 13159 9039 14244 9063
rect 11546 9033 14244 9039
rect 14480 9266 15600 9269
rect 14480 9033 14903 9266
rect 11546 9030 14903 9033
rect 15139 9235 15600 9266
rect 15836 9363 16065 9471
rect 16301 9363 16575 9599
rect 16811 9363 17084 9599
rect 17320 9363 17593 9599
rect 17829 9363 17897 9599
rect 15836 9261 17897 9363
rect 15836 9235 16065 9261
rect 15139 9139 16065 9235
rect 15139 9030 15600 9139
rect 11546 9000 15600 9030
rect 11546 8893 12226 9000
rect 10289 8837 11159 8893
rect 10013 8817 11159 8837
rect 10013 8778 10856 8817
rect 9366 8693 9625 8778
rect 8962 8550 9625 8693
rect 8605 8536 9625 8550
rect 7218 8476 8000 8536
rect 6805 8469 7132 8476
rect 4431 8432 5275 8469
rect 4431 8399 4945 8432
rect 4128 8292 4945 8399
rect 3248 8126 3746 8292
rect 0 8087 3746 8126
tri 3746 8087 3951 8292 sw
tri 4128 8087 4333 8292 ne
rect 4333 8271 4945 8292
rect 4333 8087 4556 8271
rect 0 8080 3951 8087
tri 2980 7913 3147 8080 ne
rect 3147 7913 3951 8080
tri 3951 7913 4125 8087 sw
tri 4333 7913 4507 8087 ne
rect 4507 8035 4556 8087
rect 4792 8196 4945 8271
rect 5181 8292 5275 8432
tri 5275 8292 5452 8469 sw
tri 5698 8400 5767 8469 ne
rect 5767 8400 5792 8469
tri 5792 8400 5861 8469 sw
tri 5877 8400 5946 8469 ne
rect 5946 8400 6720 8469
tri 5767 8306 5861 8400 ne
tri 5861 8391 5870 8400 sw
tri 5946 8391 5955 8400 ne
rect 5955 8391 6720 8400
rect 5861 8306 5870 8391
tri 5870 8306 5955 8391 sw
tri 5955 8306 6040 8391 ne
rect 6040 8390 6720 8391
tri 6720 8390 6799 8469 sw
tri 6805 8390 6884 8469 ne
rect 6884 8390 7132 8469
tri 7132 8390 7218 8476 sw
tri 7218 8390 7304 8476 ne
rect 7304 8451 8000 8476
tri 8000 8451 8085 8536 sw
tri 8085 8451 8170 8536 ne
rect 8170 8451 8179 8536
rect 7304 8442 8085 8451
tri 8085 8442 8094 8451 sw
tri 8170 8442 8179 8451 ne
tri 8179 8442 8273 8536 sw
tri 8605 8446 8695 8536 ne
rect 8695 8523 9625 8536
tri 9625 8523 9880 8778 sw
tri 10013 8523 10268 8778 ne
rect 10268 8674 10856 8778
rect 10268 8523 10452 8674
rect 8695 8446 9536 8523
tri 8695 8442 8699 8446 ne
rect 8699 8442 9536 8446
rect 7304 8390 8094 8442
tri 8094 8390 8146 8442 sw
tri 8179 8390 8231 8442 ne
rect 8231 8390 8273 8442
tri 8273 8390 8325 8442 sw
tri 8699 8390 8751 8442 ne
rect 8751 8390 9536 8442
rect 6040 8306 6799 8390
tri 5861 8292 5875 8306 ne
rect 5875 8297 5955 8306
tri 5955 8297 5964 8306 sw
tri 6040 8297 6049 8306 ne
rect 6049 8305 6799 8306
tri 6799 8305 6884 8390 sw
tri 6884 8305 6969 8390 ne
rect 6969 8305 7218 8390
rect 6049 8297 6884 8305
rect 5875 8292 5964 8297
tri 5964 8292 5969 8297 sw
tri 6049 8292 6054 8297 ne
rect 6054 8292 6884 8297
tri 6884 8292 6897 8305 sw
tri 6969 8292 6982 8305 ne
rect 6982 8304 7218 8305
tri 7218 8304 7304 8390 sw
tri 7304 8304 7390 8390 ne
rect 7390 8348 8146 8390
tri 8146 8348 8188 8390 sw
tri 8231 8348 8273 8390 ne
rect 8273 8348 8325 8390
tri 8325 8348 8367 8390 sw
tri 8751 8348 8793 8390 ne
rect 8793 8382 9536 8390
rect 8793 8348 9130 8382
rect 7390 8304 8188 8348
rect 6982 8292 7304 8304
tri 7304 8292 7316 8304 sw
tri 7390 8292 7402 8304 ne
rect 7402 8292 8188 8304
rect 5181 8196 5452 8292
rect 4792 8068 5452 8196
tri 5452 8068 5676 8292 sw
tri 5875 8212 5955 8292 ne
rect 5955 8212 5969 8292
tri 5969 8212 6049 8292 sw
tri 6054 8212 6134 8292 ne
rect 6134 8212 6897 8292
tri 5955 8118 6049 8212 ne
tri 6049 8203 6058 8212 sw
tri 6134 8203 6143 8212 ne
rect 6143 8207 6897 8212
tri 6897 8207 6982 8292 sw
tri 6982 8207 7067 8292 ne
rect 7067 8207 7316 8292
rect 6143 8203 6982 8207
rect 6049 8118 6058 8203
tri 6058 8118 6143 8203 sw
tri 6143 8118 6228 8203 ne
rect 6228 8141 6982 8203
tri 6982 8141 7048 8207 sw
tri 7067 8141 7133 8207 ne
rect 7133 8206 7316 8207
tri 7316 8206 7402 8292 sw
tri 7402 8206 7488 8292 ne
rect 7488 8263 8188 8292
tri 8188 8263 8273 8348 sw
tri 8273 8263 8358 8348 ne
rect 8358 8263 8367 8348
rect 7488 8254 8273 8263
tri 8273 8254 8282 8263 sw
tri 8358 8254 8367 8263 ne
tri 8367 8254 8461 8348 sw
tri 8793 8254 8887 8348 ne
rect 8887 8254 9130 8348
rect 7488 8206 8282 8254
rect 7133 8142 7402 8206
tri 7402 8142 7466 8206 sw
tri 7488 8142 7552 8206 ne
rect 7552 8169 8282 8206
tri 8282 8169 8367 8254 sw
tri 8367 8169 8452 8254 ne
rect 8452 8169 8461 8254
rect 7552 8160 8367 8169
tri 8367 8160 8376 8169 sw
tri 8452 8160 8461 8169 ne
tri 8461 8160 8555 8254 sw
tri 8887 8160 8981 8254 ne
rect 8981 8160 9130 8254
rect 7552 8142 8376 8160
rect 7133 8141 7466 8142
rect 6228 8118 7048 8141
tri 6049 8068 6099 8118 ne
rect 6099 8109 6143 8118
tri 6143 8109 6152 8118 sw
tri 6228 8109 6237 8118 ne
rect 6237 8109 7048 8118
rect 6099 8068 6152 8109
rect 4792 8035 5306 8068
rect 4507 7913 5306 8035
tri 3147 7800 3260 7913 ne
rect 3260 7831 4125 7913
tri 4125 7831 4207 7913 sw
tri 4507 7831 4589 7913 ne
rect 4589 7885 5306 7913
rect 4589 7831 4945 7885
rect 3260 7800 4207 7831
rect 0 7792 2874 7800
tri 2874 7792 2882 7800 sw
tri 3260 7792 3268 7800 ne
rect 3268 7792 4207 7800
rect 0 7738 2882 7792
rect 0 7502 277 7738
rect 513 7502 860 7738
rect 1096 7502 1442 7738
rect 1678 7502 2024 7738
rect 2260 7502 2606 7738
rect 2842 7502 2882 7738
rect 0 7496 2882 7502
tri 2882 7496 3178 7792 sw
tri 3268 7496 3564 7792 ne
rect 3564 7496 4207 7792
rect 0 7400 3178 7496
rect 0 7164 277 7400
rect 513 7164 860 7400
rect 1096 7164 1442 7400
rect 1678 7164 2024 7400
rect 2260 7164 2606 7400
rect 2842 7164 3178 7400
rect 0 7145 3178 7164
tri 3178 7145 3529 7496 sw
tri 3564 7145 3915 7496 ne
rect 3915 7449 4207 7496
tri 4207 7449 4589 7831 sw
tri 4589 7649 4771 7831 ne
rect 4771 7649 4945 7831
rect 5181 7832 5306 7885
rect 5542 7913 5676 8068
tri 5676 7913 5831 8068 sw
tri 6099 8024 6143 8068 ne
rect 6143 8024 6152 8068
tri 6152 8024 6237 8109 sw
tri 6237 8024 6322 8109 ne
rect 6322 8056 7048 8109
tri 7048 8056 7133 8141 sw
tri 7133 8056 7218 8141 ne
rect 7218 8056 7466 8141
tri 7466 8056 7552 8142 sw
tri 7552 8056 7638 8142 ne
rect 7638 8075 8376 8142
tri 8376 8075 8461 8160 sw
tri 8461 8075 8546 8160 ne
rect 8546 8075 8555 8160
rect 7638 8066 8461 8075
tri 8461 8066 8470 8075 sw
tri 8546 8066 8555 8075 ne
tri 8555 8066 8649 8160 sw
tri 8981 8146 8995 8160 ne
rect 8995 8146 9130 8160
rect 9366 8287 9536 8382
rect 9772 8506 9880 8523
tri 9880 8506 9897 8523 sw
tri 10268 8506 10285 8523 ne
rect 10285 8506 10452 8523
rect 9772 8497 9897 8506
tri 9897 8497 9906 8506 sw
tri 10285 8497 10294 8506 ne
rect 10294 8497 10452 8506
rect 9772 8390 9906 8497
tri 9906 8390 10013 8497 sw
tri 10294 8390 10401 8497 ne
rect 10401 8438 10452 8497
rect 10688 8581 10856 8674
rect 11092 8581 11159 8817
rect 10688 8506 11159 8581
tri 11159 8506 11546 8893 sw
tri 11546 8506 11933 8893 ne
rect 11933 8764 12226 8893
rect 12462 8975 15600 9000
rect 12462 8951 13547 8975
rect 12462 8764 12923 8951
rect 11933 8715 12923 8764
rect 13159 8739 13547 8951
rect 13783 8946 15600 8975
rect 13783 8739 14244 8946
rect 13159 8715 14244 8739
rect 11933 8710 14244 8715
rect 14480 8945 15600 8946
rect 14480 8710 14903 8945
rect 11933 8709 14903 8710
rect 15139 8903 15600 8945
rect 15836 9025 16065 9139
rect 16301 9025 16575 9261
rect 16811 9025 17084 9261
rect 17320 9025 17593 9261
rect 17829 9025 17897 9261
rect 15836 8923 17897 9025
rect 15836 8903 16065 8923
rect 15139 8807 16065 8903
rect 15139 8709 15600 8807
rect 11933 8675 15600 8709
rect 11933 8506 12226 8675
rect 10688 8497 11546 8506
tri 11546 8497 11555 8506 sw
tri 11933 8497 11942 8506 ne
rect 11942 8497 12226 8506
rect 10688 8438 11555 8497
rect 10401 8390 11555 8438
rect 9772 8287 10013 8390
rect 9366 8146 10013 8287
tri 8995 8066 9075 8146 ne
rect 9075 8107 10013 8146
tri 10013 8107 10296 8390 sw
tri 10401 8107 10684 8390 ne
rect 10684 8370 11555 8390
rect 10684 8270 11303 8370
rect 10684 8107 10856 8270
rect 9075 8066 9955 8107
rect 7638 8056 8470 8066
rect 6322 8024 7133 8056
tri 6143 7930 6237 8024 ne
tri 6237 8015 6246 8024 sw
tri 6322 8015 6331 8024 ne
rect 6331 8015 7133 8024
rect 6237 7930 6246 8015
tri 6246 7930 6331 8015 sw
tri 6331 7930 6416 8015 ne
rect 6416 7971 7133 8015
tri 7133 7971 7218 8056 sw
tri 7218 7971 7303 8056 ne
rect 7303 7971 7552 8056
rect 6416 7954 7218 7971
tri 7218 7954 7235 7971 sw
tri 7303 7954 7320 7971 ne
rect 7320 7970 7552 7971
tri 7552 7970 7638 8056 sw
tri 7638 7970 7724 8056 ne
rect 7724 7981 8470 8056
tri 8470 7981 8555 8066 sw
tri 8555 7981 8640 8066 ne
rect 8640 8020 8649 8066
tri 8649 8020 8695 8066 sw
tri 9075 8020 9121 8066 ne
rect 9121 8020 9955 8066
rect 8640 7981 8695 8020
rect 7724 7972 8555 7981
tri 8555 7972 8564 7981 sw
tri 8640 7972 8649 7981 ne
rect 8649 7972 8695 7981
tri 8695 7972 8743 8020 sw
tri 9121 7972 9169 8020 ne
rect 9169 7976 9955 8020
rect 9169 7972 9536 7976
rect 7724 7970 8564 7972
rect 7320 7954 7638 7970
tri 7638 7954 7654 7970 sw
tri 7724 7954 7740 7970 ne
rect 7740 7954 8564 7970
rect 6416 7930 7235 7954
tri 6237 7913 6254 7930 ne
rect 6254 7921 6331 7930
tri 6331 7921 6340 7930 sw
tri 6416 7921 6425 7930 ne
rect 6425 7926 7235 7930
tri 7235 7926 7263 7954 sw
tri 7320 7926 7348 7954 ne
rect 7348 7926 7654 7954
rect 6425 7921 7263 7926
rect 6254 7913 6340 7921
rect 5542 7832 5831 7913
rect 5181 7747 5831 7832
tri 5831 7747 5997 7913 sw
tri 6254 7836 6331 7913 ne
rect 6331 7836 6340 7913
tri 6340 7836 6425 7921 sw
tri 6425 7836 6510 7921 ne
rect 6510 7841 7263 7921
tri 7263 7841 7348 7926 sw
tri 7348 7841 7433 7926 ne
rect 7433 7868 7654 7926
tri 7654 7868 7740 7954 sw
tri 7740 7868 7826 7954 ne
rect 7826 7926 8564 7954
tri 8564 7926 8610 7972 sw
tri 8649 7926 8695 7972 ne
rect 8695 7926 8743 7972
rect 7826 7878 8610 7926
tri 8610 7878 8658 7926 sw
tri 8695 7878 8743 7926 ne
tri 8743 7878 8837 7972 sw
tri 9169 7878 9263 7972 ne
rect 9263 7878 9536 7972
rect 7826 7868 8658 7878
rect 7433 7841 7740 7868
tri 7740 7841 7767 7868 sw
tri 7826 7841 7853 7868 ne
rect 7853 7841 8658 7868
tri 8658 7841 8695 7878 sw
tri 8743 7841 8780 7878 ne
rect 8780 7841 8837 7878
tri 8837 7841 8874 7878 sw
tri 9263 7841 9300 7878 ne
rect 9300 7841 9536 7878
rect 6510 7836 7348 7841
tri 6331 7747 6420 7836 ne
rect 6420 7827 6425 7836
tri 6425 7827 6434 7836 sw
tri 6510 7827 6519 7836 ne
rect 6519 7827 7348 7836
rect 6420 7747 6434 7827
tri 6434 7747 6514 7827 sw
tri 6519 7747 6599 7827 ne
rect 6599 7807 7348 7827
tri 7348 7807 7382 7841 sw
tri 7433 7807 7467 7841 ne
rect 7467 7808 7767 7841
tri 7767 7808 7800 7841 sw
tri 7853 7808 7886 7841 ne
rect 7886 7808 8695 7841
rect 7467 7807 7800 7808
rect 6599 7747 7382 7807
rect 5181 7669 5997 7747
rect 5181 7649 5692 7669
tri 4771 7449 4971 7649 ne
rect 4971 7521 5692 7649
rect 4971 7449 5306 7521
rect 3915 7145 4589 7449
tri 4589 7145 4893 7449 sw
tri 4971 7145 5275 7449 ne
rect 5275 7285 5306 7449
rect 5542 7433 5692 7521
rect 5928 7449 5997 7669
tri 5997 7449 6295 7747 sw
tri 6420 7742 6425 7747 ne
rect 6425 7742 6514 7747
tri 6514 7742 6519 7747 sw
tri 6599 7742 6604 7747 ne
rect 6604 7742 7382 7747
tri 6425 7648 6519 7742 ne
tri 6519 7733 6528 7742 sw
tri 6604 7733 6613 7742 ne
rect 6613 7733 7382 7742
rect 6519 7648 6528 7733
tri 6528 7648 6613 7733 sw
tri 6613 7648 6698 7733 ne
rect 6698 7722 7382 7733
tri 7382 7722 7467 7807 sw
tri 7467 7722 7552 7807 ne
rect 7552 7722 7800 7807
tri 7800 7722 7886 7808 sw
tri 7886 7722 7972 7808 ne
rect 7972 7784 8695 7808
tri 8695 7784 8752 7841 sw
tri 8780 7784 8837 7841 ne
rect 8837 7784 8874 7841
tri 8874 7784 8931 7841 sw
tri 9300 7784 9357 7841 ne
rect 9357 7784 9536 7841
rect 7972 7722 8752 7784
rect 6698 7648 7467 7722
tri 6519 7554 6613 7648 ne
tri 6613 7639 6622 7648 sw
tri 6698 7639 6707 7648 ne
rect 6707 7639 7467 7648
rect 6613 7554 6622 7639
tri 6622 7554 6707 7639 sw
tri 6707 7554 6792 7639 ne
rect 6792 7637 7467 7639
tri 7467 7637 7552 7722 sw
tri 7552 7637 7637 7722 ne
rect 7637 7637 7886 7722
rect 6792 7554 7552 7637
tri 6613 7460 6707 7554 ne
tri 6707 7545 6716 7554 sw
tri 6792 7545 6801 7554 ne
rect 6801 7552 7552 7554
tri 7552 7552 7637 7637 sw
tri 7637 7552 7722 7637 ne
rect 7722 7636 7886 7637
tri 7886 7636 7972 7722 sw
tri 7972 7636 8058 7722 ne
rect 8058 7699 8752 7722
tri 8752 7699 8837 7784 sw
tri 8837 7699 8922 7784 ne
rect 8922 7699 8931 7784
rect 8058 7690 8837 7699
tri 8837 7690 8846 7699 sw
tri 8922 7690 8931 7699 ne
tri 8931 7690 9025 7784 sw
tri 9357 7740 9401 7784 ne
rect 9401 7740 9536 7784
rect 9772 7871 9955 7976
rect 10191 8002 10296 8107
tri 10296 8002 10401 8107 sw
tri 10684 8002 10789 8107 ne
rect 10789 8034 10856 8107
rect 11092 8134 11303 8270
rect 11539 8134 11555 8370
rect 11092 8110 11555 8134
tri 11555 8110 11942 8497 sw
tri 11942 8439 12000 8497 ne
rect 12000 8439 12226 8497
rect 12462 8651 15600 8675
rect 12462 8627 13547 8651
rect 12462 8439 12923 8627
tri 12000 8110 12329 8439 ne
rect 12329 8391 12923 8439
rect 13159 8415 13547 8627
rect 13783 8624 15600 8651
rect 13783 8623 14903 8624
rect 13783 8415 14244 8623
rect 13159 8391 14244 8415
rect 12329 8387 14244 8391
rect 14480 8388 14903 8623
rect 15139 8571 15600 8624
rect 15836 8687 16065 8807
rect 16301 8687 16575 8923
rect 16811 8687 17084 8923
rect 17320 8687 17593 8923
rect 17829 8687 17897 8923
rect 15836 8571 17897 8687
rect 15139 8506 17897 8571
tri 17897 8506 18991 9600 sw
rect 35157 9514 35250 9750
rect 35486 9514 35584 9750
rect 35820 9514 35918 9750
rect 36154 9514 36252 9750
rect 36488 9514 36586 9750
rect 36822 9514 36920 9750
rect 37156 9514 37254 9750
rect 37490 9514 37588 9750
rect 37824 9514 37922 9750
rect 38158 9514 38256 9750
rect 38492 9514 38590 9750
rect 38826 9514 38924 9750
rect 39160 9514 39258 9750
rect 39494 9514 39592 9750
rect 39828 9514 40000 9750
rect 35157 9428 40000 9514
rect 35157 9192 35250 9428
rect 35486 9192 35584 9428
rect 35820 9192 35918 9428
rect 36154 9192 36252 9428
rect 36488 9192 36586 9428
rect 36822 9192 36920 9428
rect 37156 9192 37254 9428
rect 37490 9192 37588 9428
rect 37824 9192 37922 9428
rect 38158 9192 38256 9428
rect 38492 9192 38590 9428
rect 38826 9192 38924 9428
rect 39160 9192 39258 9428
rect 39494 9192 39592 9428
rect 39828 9192 40000 9428
rect 35157 9106 40000 9192
rect 35157 8870 35250 9106
rect 35486 8870 35584 9106
rect 35820 8870 35918 9106
rect 36154 8870 36252 9106
rect 36488 8870 36586 9106
rect 36822 8870 36920 9106
rect 37156 8870 37254 9106
rect 37490 8870 37588 9106
rect 37824 8870 37922 9106
rect 38158 8870 38256 9106
rect 38492 8870 38590 9106
rect 38826 8870 38924 9106
rect 39160 8870 39258 9106
rect 39494 8870 39592 9106
rect 39828 8870 40000 9106
rect 35157 8784 40000 8870
rect 35157 8548 35250 8784
rect 35486 8548 35584 8784
rect 35820 8548 35918 8784
rect 36154 8548 36252 8784
rect 36488 8548 36586 8784
rect 36822 8548 36920 8784
rect 37156 8548 37254 8784
rect 37490 8548 37588 8784
rect 37824 8548 37922 8784
rect 38158 8548 38256 8784
rect 38492 8548 38590 8784
rect 38826 8548 38924 8784
rect 39160 8548 39258 8784
rect 39494 8548 39592 8784
rect 39828 8548 40000 8784
rect 15139 8501 18991 8506
rect 15139 8475 16047 8501
rect 15139 8388 15600 8475
rect 14480 8387 15600 8388
rect 12329 8327 15600 8387
rect 12329 8303 13547 8327
rect 12329 8110 12923 8303
rect 11092 8034 11942 8110
rect 10789 8019 11942 8034
tri 11942 8019 12033 8110 sw
tri 12329 8019 12420 8110 ne
rect 12420 8067 12923 8110
rect 13159 8091 13547 8303
rect 13783 8302 15600 8327
rect 13783 8300 14903 8302
rect 13783 8091 14244 8300
rect 13159 8067 14244 8091
rect 12420 8064 14244 8067
rect 14480 8066 14903 8300
rect 15139 8239 15600 8302
rect 15836 8265 16047 8475
rect 16283 8265 16549 8501
rect 16785 8265 17050 8501
rect 17286 8265 17551 8501
rect 17787 8265 18052 8501
rect 18288 8265 18553 8501
rect 18789 8497 18991 8501
tri 18991 8497 19000 8506 sw
rect 18789 8265 19000 8497
rect 15836 8239 19000 8265
rect 15139 8143 19000 8239
rect 15139 8066 15600 8143
rect 14480 8064 15600 8066
rect 12420 8019 15600 8064
rect 10789 8002 12033 8019
rect 10191 7904 10401 8002
tri 10401 7904 10499 8002 sw
tri 10789 7904 10887 8002 ne
rect 10887 7966 12033 8002
rect 10887 7904 11707 7966
rect 10191 7871 10499 7904
rect 9772 7743 10499 7871
tri 10499 7743 10660 7904 sw
tri 10887 7743 11048 7904 ne
rect 11048 7823 11707 7904
rect 11048 7743 11303 7823
rect 9772 7740 10316 7743
tri 9401 7690 9451 7740 ne
rect 9451 7690 10316 7740
rect 8058 7636 8846 7690
rect 7722 7560 7972 7636
tri 7972 7560 8048 7636 sw
tri 8058 7560 8134 7636 ne
rect 8134 7605 8846 7636
tri 8846 7605 8931 7690 sw
tri 8931 7605 9016 7690 ne
rect 9016 7605 9025 7690
rect 8134 7596 8931 7605
tri 8931 7596 8940 7605 sw
tri 9016 7596 9025 7605 ne
tri 9025 7596 9119 7690 sw
tri 9451 7604 9537 7690 ne
rect 9537 7604 10316 7690
tri 9537 7596 9545 7604 ne
rect 9545 7596 10316 7604
rect 8134 7560 8940 7596
rect 7722 7552 8048 7560
rect 6801 7545 7637 7552
rect 6707 7460 6716 7545
tri 6716 7460 6801 7545 sw
tri 6801 7460 6886 7545 ne
rect 6886 7534 7637 7545
tri 7637 7534 7655 7552 sw
tri 7722 7534 7740 7552 ne
rect 7740 7534 8048 7552
rect 6886 7460 7655 7534
tri 6707 7449 6718 7460 ne
rect 6718 7451 6801 7460
tri 6801 7451 6810 7460 sw
tri 6886 7451 6895 7460 ne
rect 6895 7451 7655 7460
rect 6718 7449 6810 7451
tri 6810 7449 6812 7451 sw
tri 6895 7449 6897 7451 ne
rect 6897 7449 7655 7451
tri 7655 7449 7740 7534 sw
tri 7740 7449 7825 7534 ne
rect 7825 7474 8048 7534
tri 8048 7474 8134 7560 sw
tri 8134 7474 8220 7560 ne
rect 8220 7511 8940 7560
tri 8940 7511 9025 7596 sw
tri 9025 7511 9110 7596 ne
rect 9110 7511 9119 7596
rect 8220 7502 9025 7511
tri 9025 7502 9034 7511 sw
tri 9110 7502 9119 7511 ne
tri 9119 7502 9213 7596 sw
tri 9545 7502 9639 7596 ne
rect 9639 7560 10316 7596
rect 9639 7502 9955 7560
rect 8220 7474 9034 7502
rect 7825 7449 8134 7474
tri 8134 7449 8159 7474 sw
tri 8220 7449 8245 7474 ne
rect 8245 7449 9034 7474
rect 5928 7433 6295 7449
rect 5542 7310 6295 7433
tri 6295 7310 6434 7449 sw
tri 6718 7366 6801 7449 ne
rect 6801 7366 6812 7449
tri 6812 7366 6895 7449 sw
tri 6897 7366 6980 7449 ne
rect 6980 7388 7740 7449
tri 7740 7388 7801 7449 sw
tri 7825 7388 7886 7449 ne
rect 7886 7388 8159 7449
tri 8159 7388 8220 7449 sw
tri 8245 7388 8306 7449 ne
rect 8306 7417 9034 7449
tri 9034 7417 9119 7502 sw
tri 9119 7417 9204 7502 ne
rect 9204 7417 9213 7502
rect 8306 7408 9119 7417
tri 9119 7408 9128 7417 sw
tri 9204 7408 9213 7417 ne
tri 9213 7408 9307 7502 sw
tri 9639 7408 9733 7502 ne
rect 9733 7408 9955 7502
rect 8306 7388 9128 7408
rect 6980 7366 7801 7388
tri 6801 7310 6857 7366 ne
rect 6857 7357 6895 7366
tri 6895 7357 6904 7366 sw
tri 6980 7357 6989 7366 ne
rect 6989 7357 7801 7366
rect 6857 7310 6904 7357
rect 5542 7285 6067 7310
rect 5275 7145 6067 7285
rect 0 7110 3529 7145
tri 3529 7110 3564 7145 sw
tri 3915 7110 3950 7145 ne
rect 3950 7110 4893 7145
tri 2588 6935 2763 7110 ne
rect 2763 6935 3564 7110
tri 3564 6935 3739 7110 sw
tri 3950 6935 4125 7110 ne
rect 4125 6935 4893 7110
tri 4893 6935 5103 7145 sw
tri 5275 6935 5485 7145 ne
rect 5485 7122 6067 7145
rect 5485 6935 5692 7122
tri 2763 6830 2868 6935 ne
rect 2868 6830 3739 6935
tri 3739 6830 3844 6935 sw
tri 4125 6830 4230 6935 ne
rect 4230 6830 5103 6935
tri 5103 6830 5208 6935 sw
tri 5485 6830 5590 6935 ne
rect 5590 6886 5692 6935
rect 5928 7074 6067 7122
rect 6303 7145 6434 7310
tri 6434 7145 6599 7310 sw
tri 6857 7272 6895 7310 ne
rect 6895 7272 6904 7310
tri 6904 7272 6989 7357 sw
tri 6989 7272 7074 7357 ne
rect 7074 7303 7801 7357
tri 7801 7303 7886 7388 sw
tri 7886 7303 7971 7388 ne
rect 7971 7303 8220 7388
rect 7074 7272 7886 7303
tri 6895 7178 6989 7272 ne
tri 6989 7263 6998 7272 sw
tri 7074 7263 7083 7272 ne
rect 7083 7263 7886 7272
rect 6989 7178 6998 7263
tri 6998 7178 7083 7263 sw
tri 7083 7178 7168 7263 ne
rect 7168 7230 7886 7263
tri 7886 7230 7959 7303 sw
tri 7971 7230 8044 7303 ne
rect 8044 7302 8220 7303
tri 8220 7302 8306 7388 sw
tri 8306 7302 8392 7388 ne
rect 8392 7323 9128 7388
tri 9128 7323 9213 7408 sw
tri 9213 7323 9298 7408 ne
rect 9298 7323 9307 7408
rect 8392 7314 9213 7323
tri 9213 7314 9222 7323 sw
tri 9298 7314 9307 7323 ne
tri 9307 7314 9401 7408 sw
tri 9733 7324 9817 7408 ne
rect 9817 7324 9955 7408
rect 10191 7507 10316 7560
rect 10552 7516 10660 7743
tri 10660 7516 10887 7743 sw
tri 11048 7516 11275 7743 ne
rect 11275 7587 11303 7743
rect 11539 7730 11707 7823
rect 11943 7730 12033 7966
rect 11539 7632 12033 7730
tri 12033 7632 12420 8019 sw
tri 12420 7632 12807 8019 ne
rect 12807 8003 15600 8019
rect 12807 7978 13547 8003
rect 12807 7742 12923 7978
rect 13159 7767 13547 7978
rect 13783 7980 15600 8003
rect 13783 7977 14903 7980
rect 13783 7767 14244 7977
rect 13159 7742 14244 7767
rect 12807 7741 14244 7742
rect 14480 7744 14903 7977
rect 15139 7907 15600 7980
rect 15836 8089 19000 8143
rect 15836 7907 16047 8089
rect 15139 7853 16047 7907
rect 16283 7853 16549 8089
rect 16785 7853 17050 8089
rect 17286 7853 17551 8089
rect 17787 7853 18052 8089
rect 18288 7853 18553 8089
rect 18789 7853 19000 8089
rect 15139 7811 19000 7853
rect 15139 7744 15600 7811
rect 14480 7741 15600 7744
rect 12807 7679 15600 7741
rect 12807 7632 13547 7679
rect 11539 7587 12420 7632
rect 11275 7567 12420 7587
rect 11275 7516 12106 7567
rect 10552 7507 10887 7516
rect 10191 7339 10887 7507
tri 10887 7339 11064 7516 sw
tri 11275 7339 11452 7516 ne
rect 11452 7419 12106 7516
rect 11452 7339 11707 7419
rect 10191 7324 10720 7339
tri 9817 7314 9827 7324 ne
rect 9827 7314 10720 7324
rect 8392 7302 9222 7314
rect 8044 7230 8306 7302
rect 7168 7178 7959 7230
tri 6989 7145 7022 7178 ne
rect 7022 7169 7083 7178
tri 7083 7169 7092 7178 sw
tri 7168 7169 7177 7178 ne
rect 7177 7169 7959 7178
rect 7022 7145 7092 7169
tri 7092 7145 7116 7169 sw
tri 7177 7145 7201 7169 ne
rect 7201 7145 7959 7169
tri 7959 7145 8044 7230 sw
tri 8044 7145 8129 7230 ne
rect 8129 7226 8306 7230
tri 8306 7226 8382 7302 sw
tri 8392 7226 8468 7302 ne
rect 8468 7229 9222 7302
tri 9222 7229 9307 7314 sw
tri 9307 7229 9392 7314 ne
rect 9392 7229 9401 7314
rect 8468 7226 9307 7229
rect 8129 7145 8382 7226
rect 6303 7074 6599 7145
rect 5928 6946 6599 7074
tri 6599 6946 6798 7145 sw
tri 7022 7084 7083 7145 ne
rect 7083 7084 7116 7145
tri 7116 7084 7177 7145 sw
tri 7201 7084 7262 7145 ne
rect 7262 7111 8044 7145
tri 8044 7111 8078 7145 sw
tri 8129 7111 8163 7145 ne
rect 8163 7140 8382 7145
tri 8382 7140 8468 7226 sw
tri 8468 7140 8554 7226 ne
rect 8554 7220 9307 7226
tri 9307 7220 9316 7229 sw
tri 9392 7220 9401 7229 ne
tri 9401 7220 9495 7314 sw
tri 9827 7220 9921 7314 ne
rect 9921 7220 10720 7314
rect 8554 7140 9316 7220
rect 8163 7111 8468 7140
tri 8468 7111 8497 7140 sw
tri 8554 7111 8583 7140 ne
rect 8583 7135 9316 7140
tri 9316 7135 9401 7220 sw
tri 9401 7135 9486 7220 ne
rect 9486 7178 9495 7220
tri 9495 7178 9537 7220 sw
tri 9921 7178 9963 7220 ne
rect 9963 7196 10720 7220
rect 9963 7178 10316 7196
rect 9486 7135 9537 7178
rect 8583 7128 9401 7135
tri 9401 7128 9408 7135 sw
tri 9486 7128 9493 7135 ne
rect 9493 7128 9537 7135
tri 9537 7128 9587 7178 sw
tri 9963 7128 10013 7178 ne
rect 10013 7128 10316 7178
rect 8583 7126 9408 7128
tri 9408 7126 9410 7128 sw
tri 9493 7126 9495 7128 ne
rect 9495 7126 9587 7128
tri 9587 7126 9589 7128 sw
tri 10013 7126 10015 7128 ne
rect 10015 7126 10316 7128
rect 8583 7111 9410 7126
rect 7262 7084 8078 7111
tri 7083 6990 7177 7084 ne
tri 7177 7075 7186 7084 sw
tri 7262 7075 7271 7084 ne
rect 7271 7075 8078 7084
rect 7177 6990 7186 7075
tri 7186 6990 7271 7075 sw
tri 7271 6990 7356 7075 ne
rect 7356 7054 8078 7075
tri 8078 7054 8135 7111 sw
tri 8163 7054 8220 7111 ne
rect 8220 7054 8497 7111
tri 8497 7054 8554 7111 sw
tri 8583 7054 8640 7111 ne
rect 8640 7084 9410 7111
tri 9410 7084 9452 7126 sw
tri 9495 7084 9537 7126 ne
rect 9537 7084 9589 7126
rect 8640 7054 9452 7084
rect 7356 6999 8135 7054
tri 8135 6999 8190 7054 sw
tri 8220 6999 8275 7054 ne
rect 8275 6999 8554 7054
tri 8554 6999 8609 7054 sw
tri 8640 6999 8695 7054 ne
rect 8695 7032 9452 7054
tri 9452 7032 9504 7084 sw
tri 9537 7032 9589 7084 ne
tri 9589 7032 9683 7126 sw
tri 10015 7032 10109 7126 ne
rect 10109 7032 10316 7126
rect 8695 6999 9504 7032
tri 9504 6999 9537 7032 sw
tri 9589 6999 9622 7032 ne
rect 9622 6999 9683 7032
tri 9683 6999 9716 7032 sw
tri 10109 6999 10142 7032 ne
rect 10142 6999 10316 7032
rect 7356 6990 8190 6999
tri 7177 6946 7221 6990 ne
rect 7221 6981 7271 6990
tri 7271 6981 7280 6990 sw
tri 7356 6981 7365 6990 ne
rect 7365 6981 8190 6990
rect 7221 6946 7280 6981
rect 5928 6886 6428 6946
rect 5590 6830 6428 6886
rect 0 6749 2472 6830
rect 0 6513 320 6749
rect 556 6513 786 6749
rect 1022 6513 1252 6749
rect 1488 6513 1718 6749
rect 1954 6513 2183 6749
rect 2419 6714 2472 6749
tri 2472 6714 2588 6830 sw
tri 2868 6714 2984 6830 ne
rect 2984 6714 3844 6830
rect 2419 6530 2588 6714
tri 2588 6530 2772 6714 sw
tri 2984 6530 3168 6714 ne
rect 3168 6530 3844 6714
rect 2419 6513 2772 6530
rect 0 6471 2772 6513
rect 0 6235 2506 6471
rect 2742 6235 2772 6471
rect 0 6215 2772 6235
rect 0 5979 320 6215
rect 556 5979 786 6215
rect 1022 5979 1252 6215
rect 1488 5979 1718 6215
rect 1954 5979 2183 6215
rect 2419 6144 2772 6215
rect 2419 5979 2506 6144
rect 0 5908 2506 5979
rect 2742 6134 2772 6144
tri 2772 6134 3168 6530 sw
tri 3168 6134 3564 6530 ne
rect 3564 6520 3844 6530
tri 3844 6520 4154 6830 sw
tri 4230 6520 4540 6830 ne
rect 4540 6763 5208 6830
tri 5208 6763 5275 6830 sw
tri 5590 6763 5657 6830 ne
rect 5657 6763 6428 6830
rect 4540 6606 5275 6763
tri 5275 6606 5432 6763 sw
tri 5657 6606 5814 6763 ne
rect 5814 6606 6067 6763
rect 4540 6520 5432 6606
rect 3564 6134 4154 6520
tri 4154 6134 4540 6520 sw
tri 4540 6134 4926 6520 ne
rect 4926 6339 5432 6520
tri 5432 6339 5699 6606 sw
tri 5814 6527 5893 6606 ne
rect 5893 6527 6067 6606
rect 6303 6710 6428 6763
rect 6664 6935 6798 6946
tri 6798 6935 6809 6946 sw
tri 7221 6935 7232 6946 ne
rect 7232 6935 7280 6946
rect 6664 6830 6809 6935
tri 6809 6830 6914 6935 sw
tri 7232 6896 7271 6935 ne
rect 7271 6896 7280 6935
tri 7280 6896 7365 6981 sw
tri 7365 6896 7450 6981 ne
rect 7450 6969 8190 6981
tri 8190 6969 8220 6999 sw
tri 8275 6969 8305 6999 ne
rect 8305 6969 8609 6999
rect 7450 6915 8220 6969
tri 8220 6915 8274 6969 sw
tri 8305 6915 8359 6969 ne
rect 8359 6915 8609 6969
rect 7450 6896 8274 6915
tri 7271 6830 7337 6896 ne
rect 7337 6887 7365 6896
tri 7365 6887 7374 6896 sw
tri 7450 6887 7459 6896 ne
rect 7459 6887 8274 6896
rect 7337 6830 7374 6887
tri 7374 6830 7431 6887 sw
tri 7459 6830 7516 6887 ne
rect 7516 6830 8274 6887
tri 8274 6830 8359 6915 sw
tri 8359 6830 8444 6915 ne
rect 8444 6913 8609 6915
tri 8609 6913 8695 6999 sw
tri 8695 6913 8781 6999 ne
rect 8781 6938 9537 6999
tri 9537 6938 9598 6999 sw
tri 9622 6938 9683 6999 ne
rect 9683 6938 9716 6999
tri 9716 6938 9777 6999 sw
tri 10142 6960 10181 6999 ne
rect 10181 6960 10316 6999
rect 10552 7103 10720 7196
rect 10956 7245 11064 7339
tri 11064 7245 11158 7339 sw
tri 11452 7245 11546 7339 ne
rect 11546 7245 11707 7339
rect 10956 7128 11158 7245
tri 11158 7128 11275 7245 sw
tri 11546 7128 11663 7245 ne
rect 11663 7183 11707 7245
rect 11943 7331 12106 7419
rect 12342 7331 12420 7567
rect 11943 7245 12420 7331
tri 12420 7245 12807 7632 sw
tri 12807 7245 13194 7632 ne
rect 13194 7443 13547 7632
rect 13783 7658 15600 7679
rect 13783 7654 14903 7658
rect 13783 7443 14244 7654
rect 13194 7418 14244 7443
rect 14480 7422 14903 7654
rect 15139 7575 15600 7658
rect 15836 7677 19000 7811
rect 15836 7575 16047 7677
rect 15139 7479 16047 7575
rect 15139 7422 15600 7479
rect 14480 7418 15600 7422
rect 13194 7354 15600 7418
rect 13194 7245 13547 7354
rect 11943 7183 12807 7245
rect 11663 7163 12807 7183
rect 11663 7128 12510 7163
rect 10956 7103 11275 7128
rect 10552 6960 11275 7103
tri 10181 6938 10203 6960 ne
rect 10203 6938 11275 6960
rect 8781 6913 9598 6938
rect 8444 6830 8695 6913
tri 8695 6830 8778 6913 sw
tri 8781 6830 8864 6913 ne
rect 8864 6853 9598 6913
tri 9598 6853 9683 6938 sw
tri 9683 6853 9768 6938 ne
rect 9768 6853 9777 6938
rect 8864 6844 9683 6853
tri 9683 6844 9692 6853 sw
tri 9768 6844 9777 6853 ne
tri 9777 6844 9871 6938 sw
tri 10203 6844 10297 6938 ne
rect 10297 6933 11275 6938
tri 11275 6933 11470 7128 sw
tri 11663 6933 11858 7128 ne
rect 11858 7020 12510 7128
rect 11858 6933 12106 7020
rect 10297 6844 11126 6933
rect 8864 6830 9692 6844
tri 9692 6830 9706 6844 sw
tri 9777 6830 9791 6844 ne
rect 9791 6830 9871 6844
rect 6664 6710 6914 6830
rect 6303 6606 6914 6710
tri 6914 6606 7138 6830 sw
tri 7337 6802 7365 6830 ne
rect 7365 6802 7431 6830
tri 7431 6802 7459 6830 sw
tri 7516 6802 7544 6830 ne
rect 7544 6805 8359 6830
tri 8359 6805 8384 6830 sw
tri 8444 6805 8469 6830 ne
rect 8469 6806 8778 6830
tri 8778 6806 8802 6830 sw
tri 8864 6806 8888 6830 ne
rect 8888 6806 9706 6830
rect 8469 6805 8802 6806
rect 7544 6802 8384 6805
tri 7365 6708 7459 6802 ne
tri 7459 6793 7468 6802 sw
tri 7544 6793 7553 6802 ne
rect 7553 6793 8384 6802
rect 7459 6708 7468 6793
tri 7468 6708 7553 6793 sw
tri 7553 6708 7638 6793 ne
rect 7638 6720 8384 6793
tri 8384 6720 8469 6805 sw
tri 8469 6720 8554 6805 ne
rect 8554 6720 8802 6805
tri 8802 6720 8888 6806 sw
tri 8888 6720 8974 6806 ne
rect 8974 6750 9706 6806
tri 9706 6750 9786 6830 sw
tri 9791 6750 9871 6830 ne
tri 9871 6750 9965 6844 sw
tri 10297 6762 10379 6844 ne
rect 10379 6792 11126 6844
rect 10379 6762 10720 6792
tri 10379 6750 10391 6762 ne
rect 10391 6750 10720 6762
rect 8974 6720 9786 6750
rect 7638 6708 8469 6720
tri 7459 6614 7553 6708 ne
tri 7553 6699 7562 6708 sw
tri 7638 6699 7647 6708 ne
rect 7647 6699 8469 6708
rect 7553 6614 7562 6699
tri 7562 6614 7647 6699 sw
tri 7647 6614 7732 6699 ne
rect 7732 6635 8469 6699
tri 8469 6635 8554 6720 sw
tri 8554 6635 8639 6720 ne
rect 8639 6635 8888 6720
rect 7732 6614 8554 6635
tri 7553 6606 7561 6614 ne
rect 7561 6606 7647 6614
tri 7647 6606 7655 6614 sw
tri 7732 6606 7740 6614 ne
rect 7740 6606 8554 6614
tri 8554 6606 8583 6635 sw
tri 8639 6606 8668 6635 ne
rect 8668 6634 8888 6635
tri 8888 6634 8974 6720 sw
tri 8974 6634 9060 6720 ne
rect 9060 6665 9786 6720
tri 9786 6665 9871 6750 sw
tri 9871 6665 9956 6750 ne
rect 9956 6665 9965 6750
rect 9060 6656 9871 6665
tri 9871 6656 9880 6665 sw
tri 9956 6656 9965 6665 ne
tri 9965 6656 10059 6750 sw
tri 10391 6656 10485 6750 ne
rect 10485 6656 10720 6750
rect 9060 6634 9880 6656
rect 8668 6606 8974 6634
tri 8974 6606 9002 6634 sw
tri 9060 6606 9088 6634 ne
rect 9088 6606 9880 6634
rect 6303 6560 7138 6606
rect 6303 6527 6817 6560
tri 5893 6339 6081 6527 ne
rect 6081 6399 6817 6527
rect 6081 6339 6428 6399
rect 4926 6134 5699 6339
rect 2742 6089 3168 6134
rect 2742 5908 2888 6089
rect 0 5900 2888 5908
tri 2075 5866 2109 5900 ne
rect 2109 5866 2888 5900
tri 2109 5620 2355 5866 ne
rect 2355 5853 2888 5866
rect 3124 5900 3168 6089
tri 3168 5900 3402 6134 sw
tri 3564 5957 3741 6134 ne
rect 3741 5957 4540 6134
tri 4540 5957 4717 6134 sw
tri 4926 5957 5103 6134 ne
rect 5103 5957 5699 6134
tri 5699 5957 6081 6339 sw
tri 6081 6163 6257 6339 ne
rect 6257 6163 6428 6339
rect 6664 6324 6817 6399
rect 7053 6423 7138 6560
tri 7138 6423 7321 6606 sw
tri 7561 6520 7647 6606 ne
rect 7647 6605 7655 6606
tri 7655 6605 7656 6606 sw
tri 7740 6605 7741 6606 ne
rect 7741 6605 8583 6606
rect 7647 6520 7656 6605
tri 7656 6520 7741 6605 sw
tri 7741 6520 7826 6605 ne
rect 7826 6521 8583 6605
tri 8583 6521 8668 6606 sw
tri 8668 6521 8753 6606 ne
rect 8753 6521 9002 6606
rect 7826 6520 8668 6521
tri 7647 6426 7741 6520 ne
tri 7741 6511 7750 6520 sw
tri 7826 6511 7835 6520 ne
rect 7835 6511 8668 6520
rect 7741 6426 7750 6511
tri 7750 6426 7835 6511 sw
tri 7835 6426 7920 6511 ne
rect 7920 6471 8668 6511
tri 8668 6471 8718 6521 sw
tri 8753 6471 8803 6521 ne
rect 8803 6520 9002 6521
tri 9002 6520 9088 6606 sw
tri 9088 6520 9174 6606 ne
rect 9174 6571 9880 6606
tri 9880 6571 9965 6656 sw
tri 9965 6571 10050 6656 ne
rect 10050 6571 10059 6656
rect 9174 6562 9965 6571
tri 9965 6562 9974 6571 sw
tri 10050 6562 10059 6571 ne
tri 10059 6562 10153 6656 sw
tri 10485 6562 10579 6656 ne
rect 10579 6562 10720 6656
rect 9174 6520 9974 6562
rect 8803 6472 9088 6520
tri 9088 6472 9136 6520 sw
tri 9174 6472 9222 6520 ne
rect 9222 6477 9974 6520
tri 9974 6477 10059 6562 sw
tri 10059 6477 10144 6562 ne
rect 10144 6477 10153 6562
rect 9222 6472 10059 6477
rect 8803 6471 9136 6472
rect 7920 6426 8718 6471
tri 7741 6423 7744 6426 ne
rect 7744 6423 7835 6426
tri 7835 6423 7838 6426 sw
tri 7920 6423 7923 6426 ne
rect 7923 6423 8718 6426
rect 7053 6332 7321 6423
tri 7321 6332 7412 6423 sw
tri 7744 6332 7835 6423 ne
rect 7835 6417 7838 6423
tri 7838 6417 7844 6423 sw
tri 7923 6417 7929 6423 ne
rect 7929 6417 8718 6423
rect 7835 6332 7844 6417
tri 7844 6332 7929 6417 sw
tri 7929 6332 8014 6417 ne
rect 8014 6386 8718 6417
tri 8718 6386 8803 6471 sw
tri 8803 6386 8888 6471 ne
rect 8888 6386 9136 6471
tri 9136 6386 9222 6472 sw
tri 9222 6386 9308 6472 ne
rect 9308 6468 10059 6472
tri 10059 6468 10068 6477 sw
tri 10144 6468 10153 6477 ne
tri 10153 6468 10247 6562 sw
tri 10579 6556 10585 6562 ne
rect 10585 6556 10720 6562
rect 10956 6697 11126 6792
rect 11362 6740 11470 6933
tri 11470 6740 11663 6933 sw
tri 11858 6740 12051 6933 ne
rect 12051 6784 12106 6933
rect 12342 6927 12510 7020
rect 12746 6927 12807 7163
rect 12342 6858 12807 6927
tri 12807 6858 13194 7245 sw
tri 13194 7118 13321 7245 ne
rect 13321 7118 13547 7245
rect 13783 7336 15600 7354
rect 13783 7331 14903 7336
rect 13783 7118 14244 7331
tri 13321 6858 13581 7118 ne
rect 13581 7095 14244 7118
rect 14480 7100 14903 7331
rect 15139 7243 15600 7336
rect 15836 7441 16047 7479
rect 16283 7441 16549 7677
rect 16785 7441 17050 7677
rect 17286 7441 17551 7677
rect 17787 7441 18052 7677
rect 18288 7441 18553 7677
rect 18789 7441 19000 7677
rect 15836 7265 19000 7441
rect 15836 7243 16047 7265
rect 15139 7147 16047 7243
rect 15139 7100 15600 7147
rect 14480 7095 15600 7100
rect 13581 6911 15600 7095
rect 15836 7029 16047 7147
rect 16283 7029 16549 7265
rect 16785 7029 17050 7265
rect 17286 7029 17551 7265
rect 17787 7029 18052 7265
rect 18288 7029 18553 7265
rect 18789 7029 19000 7265
rect 15836 6911 19000 7029
rect 13581 6858 19000 6911
rect 12342 6784 13194 6858
rect 12051 6740 13194 6784
rect 11362 6697 11663 6740
rect 10956 6556 11663 6697
tri 10585 6468 10673 6556 ne
rect 10673 6468 11663 6556
rect 9308 6386 10068 6468
rect 8014 6332 8803 6386
rect 7053 6324 7412 6332
rect 6664 6196 7412 6324
tri 7412 6196 7548 6332 sw
tri 7835 6238 7929 6332 ne
tri 7929 6323 7938 6332 sw
tri 8014 6323 8023 6332 ne
rect 8023 6323 8803 6332
rect 7929 6238 7938 6323
tri 7938 6238 8023 6323 sw
tri 8023 6238 8108 6323 ne
rect 8108 6301 8803 6323
tri 8803 6301 8888 6386 sw
tri 8888 6301 8973 6386 ne
rect 8973 6301 9222 6386
rect 8108 6268 8888 6301
tri 8888 6268 8921 6301 sw
tri 8973 6268 9006 6301 ne
rect 9006 6300 9222 6301
tri 9222 6300 9308 6386 sw
tri 9308 6300 9394 6386 ne
rect 9394 6383 10068 6386
tri 10068 6383 10153 6468 sw
tri 10153 6383 10238 6468 ne
rect 10238 6383 10247 6468
rect 9394 6374 10153 6383
tri 10153 6374 10162 6383 sw
tri 10238 6374 10247 6383 ne
tri 10247 6374 10341 6468 sw
tri 10673 6374 10767 6468 ne
rect 10767 6432 11663 6468
tri 11663 6432 11971 6740 sw
tri 12051 6432 12359 6740 ne
rect 12359 6732 13194 6740
tri 13194 6732 13320 6858 sw
tri 13581 6732 13707 6858 ne
rect 13707 6853 19000 6858
rect 13707 6732 16047 6853
rect 12359 6616 13320 6732
rect 12359 6432 12510 6616
rect 10767 6386 11971 6432
rect 10767 6374 11126 6386
rect 9394 6300 10162 6374
rect 9006 6268 9308 6300
tri 9308 6268 9340 6300 sw
tri 9394 6268 9426 6300 ne
rect 9426 6289 10162 6300
tri 10162 6289 10247 6374 sw
tri 10247 6289 10332 6374 ne
rect 10332 6336 10341 6374
tri 10341 6336 10379 6374 sw
tri 10767 6336 10805 6374 ne
rect 10805 6336 11126 6374
rect 10332 6289 10379 6336
rect 9426 6280 10247 6289
tri 10247 6280 10256 6289 sw
tri 10332 6280 10341 6289 ne
rect 10341 6280 10379 6289
tri 10379 6280 10435 6336 sw
tri 10805 6280 10861 6336 ne
rect 10861 6280 11126 6336
rect 9426 6268 10256 6280
rect 8108 6242 8921 6268
tri 8921 6242 8947 6268 sw
tri 9006 6242 9032 6268 ne
rect 9032 6242 9340 6268
rect 8108 6238 8947 6242
tri 7929 6196 7971 6238 ne
rect 7971 6229 8023 6238
tri 8023 6229 8032 6238 sw
tri 8108 6229 8117 6238 ne
rect 8117 6229 8947 6238
rect 7971 6196 8032 6229
rect 6664 6163 7178 6196
tri 6257 5957 6463 6163 ne
rect 6463 6013 7178 6163
rect 6463 5957 6817 6013
tri 3741 5900 3798 5957 ne
rect 3798 5900 4717 5957
tri 4717 5900 4774 5957 sw
tri 5103 5900 5160 5957 ne
rect 5160 5900 6081 5957
tri 6081 5900 6138 5957 sw
tri 6463 5900 6520 5957 ne
rect 6520 5900 6817 5957
rect 3124 5866 3402 5900
tri 3402 5866 3436 5900 sw
tri 3798 5866 3832 5900 ne
rect 3832 5866 4774 5900
tri 4774 5866 4808 5900 sw
tri 5160 5866 5194 5900 ne
rect 5194 5866 6138 5900
tri 6138 5866 6172 5900 sw
tri 6520 5866 6554 5900 ne
rect 6554 5866 6817 5900
rect 3124 5853 3436 5866
rect 2355 5816 3436 5853
rect 2355 5620 2506 5816
rect 0 5542 1961 5620
rect 0 5306 305 5542
rect 541 5306 772 5542
rect 1008 5306 1239 5542
rect 1475 5306 1706 5542
rect 1942 5494 1961 5542
tri 1961 5494 2087 5620 sw
tri 2355 5494 2481 5620 ne
rect 2481 5580 2506 5620
rect 2742 5762 3436 5816
rect 2742 5580 2888 5762
rect 2481 5526 2888 5580
rect 3124 5738 3436 5762
tri 3436 5738 3564 5866 sw
tri 3832 5821 3877 5866 ne
rect 3877 5821 4808 5866
tri 4808 5821 4853 5866 sw
tri 5194 5821 5239 5866 ne
rect 5239 5821 6172 5866
tri 6172 5821 6217 5866 sw
tri 6554 5821 6599 5866 ne
rect 6599 5821 6817 5866
tri 3877 5738 3960 5821 ne
rect 3960 5738 4853 5821
rect 3124 5676 3564 5738
rect 3124 5526 3301 5676
rect 2481 5494 3301 5526
rect 1942 5306 2087 5494
rect 0 5121 2087 5306
tri 2087 5121 2460 5494 sw
tri 2481 5121 2854 5494 ne
rect 2854 5440 3301 5494
rect 3537 5494 3564 5676
tri 3564 5494 3808 5738 sw
tri 3960 5494 4204 5738 ne
rect 4204 5544 4853 5738
tri 4853 5544 5130 5821 sw
tri 5239 5544 5516 5821 ne
rect 5516 5763 6217 5821
tri 6217 5763 6275 5821 sw
tri 6599 5763 6657 5821 ne
rect 6657 5777 6817 5821
rect 7053 5960 7178 6013
rect 7414 5960 7548 6196
rect 7053 5957 7548 5960
tri 7548 5957 7787 6196 sw
tri 7971 6144 8023 6196 ne
rect 8023 6144 8032 6196
tri 8032 6144 8117 6229 sw
tri 8117 6144 8202 6229 ne
rect 8202 6157 8947 6229
tri 8947 6157 9032 6242 sw
tri 9032 6157 9117 6242 ne
rect 9117 6182 9340 6242
tri 9340 6182 9426 6268 sw
tri 9426 6182 9512 6268 ne
rect 9512 6242 10256 6268
tri 10256 6242 10294 6280 sw
tri 10341 6242 10379 6280 ne
rect 10379 6242 10435 6280
rect 9512 6186 10294 6242
tri 10294 6186 10350 6242 sw
tri 10379 6186 10435 6242 ne
tri 10435 6186 10529 6280 sw
tri 10861 6186 10955 6280 ne
rect 10955 6186 11126 6280
rect 9512 6182 10350 6186
rect 9117 6157 9426 6182
tri 9426 6157 9451 6182 sw
tri 9512 6157 9537 6182 ne
rect 9537 6157 10350 6182
tri 10350 6157 10379 6186 sw
tri 10435 6157 10464 6186 ne
rect 10464 6157 10529 6186
tri 10529 6157 10558 6186 sw
tri 10955 6157 10984 6186 ne
rect 10984 6157 11126 6186
rect 8202 6144 9032 6157
tri 8023 6050 8117 6144 ne
tri 8117 6135 8126 6144 sw
tri 8202 6135 8211 6144 ne
rect 8211 6137 9032 6144
tri 9032 6137 9052 6157 sw
tri 9117 6137 9137 6157 ne
rect 9137 6138 9451 6157
tri 9451 6138 9470 6157 sw
tri 9537 6138 9556 6157 ne
rect 9556 6138 10379 6157
rect 9137 6137 9470 6138
rect 8211 6135 9052 6137
rect 8117 6050 8126 6135
tri 8126 6050 8211 6135 sw
tri 8211 6050 8296 6135 ne
rect 8296 6052 9052 6135
tri 9052 6052 9137 6137 sw
tri 9137 6052 9222 6137 ne
rect 9222 6052 9470 6137
tri 9470 6052 9556 6138 sw
tri 9556 6052 9642 6138 ne
rect 9642 6092 10379 6138
tri 10379 6092 10444 6157 sw
tri 10464 6092 10529 6157 ne
rect 10529 6092 10558 6157
tri 10558 6092 10623 6157 sw
tri 10984 6150 10991 6157 ne
rect 10991 6150 11126 6157
rect 11362 6254 11971 6386
tri 11971 6254 12149 6432 sw
tri 12359 6380 12411 6432 ne
rect 12411 6380 12510 6432
rect 12746 6432 13320 6616
tri 13320 6432 13620 6732 sw
tri 13707 6432 14007 6732 ne
rect 14007 6617 16047 6732
rect 16283 6617 16549 6853
rect 16785 6617 17050 6853
rect 17286 6617 17551 6853
rect 17787 6617 18052 6853
rect 18288 6617 18553 6853
rect 18789 6617 19000 6853
rect 14007 6489 19000 6617
rect 12746 6380 13620 6432
tri 12411 6254 12537 6380 ne
rect 12537 6345 13620 6380
tri 13620 6345 13707 6432 sw
rect 12537 6279 13707 6345
rect 12537 6254 12869 6279
rect 11362 6150 12149 6254
tri 10991 6092 11049 6150 ne
rect 11049 6092 12149 6150
rect 9642 6052 10444 6092
rect 8296 6050 9137 6052
tri 8117 5957 8210 6050 ne
rect 8210 6041 8211 6050
tri 8211 6041 8220 6050 sw
tri 8296 6041 8305 6050 ne
rect 8305 6041 9137 6050
rect 8210 5957 8220 6041
rect 7053 5900 7787 5957
tri 7787 5900 7844 5957 sw
tri 8210 5956 8211 5957 ne
rect 8211 5956 8220 5957
tri 8220 5956 8305 6041 sw
tri 8305 5956 8390 6041 ne
rect 8390 5967 9137 6041
tri 9137 5967 9222 6052 sw
tri 9222 5967 9307 6052 ne
rect 9307 5967 9556 6052
rect 8390 5956 9222 5967
tri 8211 5900 8267 5956 ne
rect 8267 5947 8305 5956
tri 8305 5947 8314 5956 sw
tri 8390 5947 8399 5956 ne
rect 8399 5947 9222 5956
rect 8267 5900 8314 5947
tri 8314 5900 8361 5947 sw
tri 8399 5900 8446 5947 ne
rect 8446 5900 9222 5947
tri 9222 5900 9289 5967 sw
tri 9307 5900 9374 5967 ne
rect 9374 5966 9556 5967
tri 9556 5966 9642 6052 sw
tri 9642 5966 9728 6052 ne
rect 9728 6007 10444 6052
tri 10444 6007 10529 6092 sw
tri 10529 6007 10614 6092 ne
rect 10614 6007 10623 6092
rect 9728 5998 10529 6007
tri 10529 5998 10538 6007 sw
tri 10614 5998 10623 6007 ne
tri 10623 5998 10717 6092 sw
tri 11049 5998 11143 6092 ne
rect 11143 5998 12149 6092
rect 9728 5966 10538 5998
rect 9374 5900 9642 5966
tri 9642 5900 9708 5966 sw
tri 9728 5900 9794 5966 ne
rect 9794 5913 10538 5966
tri 10538 5913 10623 5998 sw
tri 10623 5913 10708 5998 ne
rect 10708 5913 10717 5998
rect 9794 5904 10623 5913
tri 10623 5904 10632 5913 sw
tri 10708 5904 10717 5913 ne
tri 10717 5904 10811 5998 sw
tri 11143 5920 11221 5998 ne
rect 11221 5984 12149 5998
tri 12149 5984 12419 6254 sw
tri 12537 5984 12807 6254 ne
rect 12807 6043 12869 6254
rect 13105 6043 13421 6279
rect 13657 6043 13707 6279
rect 12807 5984 13707 6043
rect 11221 5974 12419 5984
tri 12419 5974 12429 5984 sw
tri 12807 5974 12817 5984 ne
rect 11221 5920 12429 5974
tri 11221 5904 11237 5920 ne
rect 11237 5904 12429 5920
rect 9794 5900 10632 5904
tri 10632 5900 10636 5904 sw
tri 10717 5900 10721 5904 ne
rect 10721 5900 10811 5904
rect 7053 5866 7844 5900
tri 7844 5866 7878 5900 sw
tri 8267 5866 8301 5900 ne
rect 8301 5866 8361 5900
tri 8361 5866 8395 5900 sw
tri 8446 5866 8480 5900 ne
rect 8480 5866 9289 5900
tri 9289 5866 9323 5900 sw
tri 9374 5866 9408 5900 ne
rect 9408 5866 9708 5900
tri 9708 5866 9742 5900 sw
tri 9794 5866 9828 5900 ne
rect 9828 5866 10636 5900
tri 10636 5866 10670 5900 sw
tri 10721 5866 10755 5900 ne
rect 10755 5866 10811 5900
tri 10811 5866 10849 5904 sw
tri 11237 5866 11275 5904 ne
rect 11275 5866 12429 5904
tri 12429 5866 12537 5974 sw
rect 7053 5821 7878 5866
tri 7878 5821 7923 5866 sw
tri 8301 5862 8305 5866 ne
rect 8305 5862 8395 5866
tri 8395 5862 8399 5866 sw
tri 8480 5862 8484 5866 ne
rect 8484 5862 9323 5866
tri 8305 5821 8346 5862 ne
rect 8346 5853 8399 5862
tri 8399 5853 8408 5862 sw
tri 8484 5853 8493 5862 ne
rect 8493 5853 9323 5862
rect 8346 5821 8408 5853
tri 8408 5821 8440 5853 sw
tri 8493 5821 8525 5853 ne
rect 8525 5848 9323 5853
tri 9323 5848 9341 5866 sw
tri 9408 5848 9426 5866 ne
rect 9426 5848 9742 5866
rect 8525 5821 9341 5848
rect 7053 5788 7923 5821
rect 7053 5777 7589 5788
rect 6657 5763 7589 5777
rect 5516 5544 6275 5763
rect 4204 5494 5130 5544
tri 5130 5494 5180 5544 sw
tri 5516 5494 5566 5544 ne
rect 5566 5494 6275 5544
tri 6275 5494 6544 5763 sw
tri 6657 5494 6926 5763 ne
rect 6926 5649 7589 5763
rect 6926 5494 7178 5649
rect 3537 5440 3808 5494
rect 2854 5434 3808 5440
rect 2854 5198 2888 5434
rect 3124 5349 3808 5434
rect 3124 5198 3301 5349
rect 2854 5121 3301 5198
rect 0 4980 2139 5121
rect 0 4744 305 4980
rect 541 4744 772 4980
rect 1008 4744 1239 4980
rect 1475 4744 1706 4980
rect 1942 4885 2139 4980
rect 2375 5100 2460 5121
tri 2460 5100 2481 5121 sw
tri 2854 5100 2875 5121 ne
rect 2875 5113 3301 5121
rect 3537 5294 3808 5349
tri 3808 5294 4008 5494 sw
tri 4204 5294 4404 5494 ne
rect 4404 5294 5180 5494
rect 3537 5113 3683 5294
rect 2875 5100 3683 5113
rect 2375 5084 2481 5100
tri 2481 5084 2497 5100 sw
tri 2875 5084 2891 5100 ne
rect 2891 5084 3683 5100
rect 2375 4885 2497 5084
rect 1942 4794 2497 4885
rect 1942 4744 2139 4794
rect 0 4690 2139 4744
tri 1584 4573 1701 4690 ne
rect 1701 4573 2139 4690
tri 1701 4410 1864 4573 ne
rect 1864 4558 2139 4573
rect 2375 4739 2497 4794
tri 2497 4739 2842 5084 sw
tri 2891 4739 3236 5084 ne
rect 3236 5058 3683 5084
rect 3919 5158 4008 5294
tri 4008 5158 4144 5294 sw
tri 4404 5158 4540 5294 ne
rect 4540 5158 5180 5294
tri 5180 5158 5516 5494 sw
tri 5566 5158 5902 5494 ne
rect 5902 5439 6544 5494
tri 6544 5439 6599 5494 sw
tri 6926 5439 6981 5494 ne
rect 6981 5439 7178 5494
rect 5902 5361 6599 5439
tri 6599 5361 6677 5439 sw
tri 6981 5361 7059 5439 ne
rect 7059 5413 7178 5439
rect 7414 5552 7589 5649
rect 7825 5763 7923 5788
tri 7923 5763 7981 5821 sw
tri 8346 5768 8399 5821 ne
rect 8399 5768 8440 5821
tri 8440 5768 8493 5821 sw
tri 8525 5768 8578 5821 ne
rect 8578 5768 9341 5821
tri 8399 5763 8404 5768 ne
rect 8404 5763 8493 5768
tri 8493 5763 8498 5768 sw
tri 8578 5763 8583 5768 ne
rect 8583 5763 9341 5768
tri 9341 5763 9426 5848 sw
tri 9426 5763 9511 5848 ne
rect 9511 5804 9742 5848
tri 9742 5804 9804 5866 sw
tri 9828 5804 9890 5866 ne
rect 9890 5810 10670 5866
tri 10670 5810 10726 5866 sw
tri 10755 5810 10811 5866 ne
rect 10811 5810 10849 5866
tri 10849 5810 10905 5866 sw
tri 11275 5810 11331 5866 ne
rect 11331 5812 12537 5866
rect 11331 5810 11703 5812
rect 9890 5804 10726 5810
rect 9511 5763 9804 5804
tri 9804 5763 9845 5804 sw
tri 9890 5763 9931 5804 ne
rect 9931 5763 10726 5804
rect 7825 5552 7981 5763
rect 7414 5494 7981 5552
tri 7981 5494 8250 5763 sw
tri 8404 5674 8493 5763 ne
rect 8493 5759 8498 5763
tri 8498 5759 8502 5763 sw
tri 8583 5759 8587 5763 ne
rect 8587 5759 9426 5763
rect 8493 5674 8502 5759
tri 8502 5674 8587 5759 sw
tri 8587 5674 8672 5759 ne
rect 8672 5718 9426 5759
tri 9426 5718 9471 5763 sw
tri 9511 5718 9556 5763 ne
rect 9556 5718 9845 5763
tri 9845 5718 9890 5763 sw
tri 9931 5718 9976 5763 ne
rect 9976 5725 10726 5763
tri 10726 5725 10811 5810 sw
tri 10811 5725 10896 5810 ne
rect 10896 5725 10905 5810
rect 9976 5718 10811 5725
rect 8672 5674 9471 5718
tri 8493 5580 8587 5674 ne
tri 8587 5665 8596 5674 sw
tri 8672 5665 8681 5674 ne
rect 8681 5665 9471 5674
rect 8587 5580 8596 5665
tri 8596 5580 8681 5665 sw
tri 8681 5580 8766 5665 ne
rect 8766 5633 9471 5665
tri 9471 5633 9556 5718 sw
tri 9556 5633 9641 5718 ne
rect 9641 5633 9890 5718
rect 8766 5580 9556 5633
tri 8587 5494 8673 5580 ne
rect 8673 5571 8681 5580
tri 8681 5571 8690 5580 sw
tri 8766 5571 8775 5580 ne
rect 8775 5579 9556 5580
tri 9556 5579 9610 5633 sw
tri 9641 5579 9695 5633 ne
rect 9695 5632 9890 5633
tri 9890 5632 9976 5718 sw
tri 9976 5632 10062 5718 ne
rect 10062 5716 10811 5718
tri 10811 5716 10820 5725 sw
tri 10896 5716 10905 5725 ne
tri 10905 5716 10999 5810 sw
tri 11331 5716 11425 5810 ne
rect 11425 5716 11703 5810
rect 10062 5632 10820 5716
rect 9695 5580 9976 5632
tri 9976 5580 10028 5632 sw
tri 10062 5580 10114 5632 ne
rect 10114 5631 10820 5632
tri 10820 5631 10905 5716 sw
tri 10905 5631 10990 5716 ne
rect 10990 5631 10999 5716
rect 10114 5622 10905 5631
tri 10905 5622 10914 5631 sw
tri 10990 5622 10999 5631 ne
tri 10999 5622 11093 5716 sw
tri 11425 5622 11519 5716 ne
rect 11519 5622 11703 5716
rect 10114 5580 10914 5622
rect 9695 5579 10028 5580
rect 8775 5571 9610 5579
rect 8673 5494 8690 5571
tri 8690 5494 8767 5571 sw
tri 8775 5494 8852 5571 ne
rect 8852 5494 9610 5571
tri 9610 5494 9695 5579 sw
tri 9695 5494 9780 5579 ne
rect 9780 5494 10028 5579
tri 10028 5494 10114 5580 sw
tri 10114 5494 10200 5580 ne
rect 10200 5537 10914 5580
tri 10914 5537 10999 5622 sw
tri 10999 5537 11084 5622 ne
rect 11084 5537 11093 5622
rect 10200 5528 10999 5537
tri 10999 5528 11008 5537 sw
tri 11084 5528 11093 5537 ne
tri 11093 5528 11187 5622 sw
tri 11519 5528 11613 5622 ne
rect 11613 5576 11703 5622
rect 11939 5576 12237 5812
rect 12473 5576 12537 5812
rect 11613 5528 12537 5576
rect 10200 5494 11008 5528
tri 11008 5494 11042 5528 sw
tri 11093 5494 11127 5528 ne
rect 11127 5494 11187 5528
tri 11187 5494 11221 5528 sw
tri 11613 5494 11647 5528 ne
rect 7414 5486 8250 5494
tri 8250 5486 8258 5494 sw
tri 8673 5486 8681 5494 ne
rect 8681 5486 8767 5494
tri 8767 5486 8775 5494 sw
tri 8852 5486 8860 5494 ne
rect 8860 5486 9695 5494
rect 7414 5424 8258 5486
rect 7414 5413 7950 5424
rect 7059 5361 7950 5413
rect 5902 5158 6677 5361
rect 3919 5058 4144 5158
rect 3236 5021 4144 5058
rect 3236 4785 3301 5021
rect 3537 4967 4144 5021
rect 3537 4785 3683 4967
rect 3236 4739 3683 4785
rect 2375 4558 2521 4739
rect 1864 4503 2521 4558
rect 2757 4690 2842 4739
tri 2842 4690 2891 4739 sw
tri 3236 4690 3285 4739 ne
rect 3285 4731 3683 4739
rect 3919 4846 4144 4967
tri 4144 4846 4456 5158 sw
tri 4540 4979 4719 5158 ne
rect 4719 4979 5516 5158
tri 5516 4979 5695 5158 sw
tri 5902 4979 6081 5158 ne
rect 6081 4979 6677 5158
tri 6677 4979 7059 5361 sw
tri 7059 4979 7441 5361 ne
rect 7441 5241 7950 5361
rect 7441 5005 7589 5241
rect 7825 5188 7950 5241
rect 8186 5188 8258 5424
rect 7825 5099 8258 5188
tri 8258 5099 8645 5486 sw
tri 8681 5392 8775 5486 ne
tri 8775 5477 8784 5486 sw
tri 8860 5477 8869 5486 ne
rect 8869 5477 9695 5486
rect 8775 5392 8784 5477
tri 8784 5392 8869 5477 sw
tri 8869 5392 8954 5477 ne
rect 8954 5425 9695 5477
tri 9695 5425 9764 5494 sw
tri 9780 5425 9849 5494 ne
rect 9849 5470 10114 5494
tri 10114 5470 10138 5494 sw
tri 10200 5470 10224 5494 ne
rect 10224 5470 11042 5494
rect 9849 5425 10138 5470
tri 10138 5425 10183 5470 sw
tri 10224 5425 10269 5470 ne
rect 10269 5434 11042 5470
tri 11042 5434 11102 5494 sw
tri 11127 5434 11187 5494 ne
rect 11187 5434 11221 5494
tri 11221 5434 11281 5494 sw
rect 11647 5487 12537 5528
rect 10269 5425 11102 5434
rect 8954 5392 9764 5425
tri 8775 5298 8869 5392 ne
tri 8869 5383 8878 5392 sw
tri 8954 5383 8963 5392 ne
rect 8963 5384 9764 5392
tri 9764 5384 9805 5425 sw
tri 9849 5384 9890 5425 ne
rect 9890 5384 10183 5425
tri 10183 5384 10224 5425 sw
tri 10269 5384 10310 5425 ne
rect 10310 5400 11102 5425
tri 11102 5400 11136 5434 sw
tri 11187 5400 11221 5434 ne
rect 11221 5400 11281 5434
rect 10310 5384 11136 5400
rect 8963 5383 9805 5384
rect 8869 5298 8878 5383
tri 8878 5298 8963 5383 sw
tri 8963 5298 9048 5383 ne
rect 9048 5315 9805 5383
tri 9805 5315 9874 5384 sw
tri 9890 5315 9959 5384 ne
rect 9959 5365 10224 5384
tri 10224 5365 10243 5384 sw
tri 10310 5365 10329 5384 ne
rect 10329 5365 11136 5384
rect 9959 5315 10243 5365
tri 10243 5315 10293 5365 sw
tri 10329 5315 10379 5365 ne
rect 10379 5340 11136 5365
tri 11136 5340 11196 5400 sw
tri 11221 5340 11281 5400 ne
tri 11281 5368 11347 5434 sw
rect 10379 5315 11196 5340
tri 11196 5315 11221 5340 sw
rect 9048 5299 9874 5315
tri 9874 5299 9890 5315 sw
tri 9959 5299 9975 5315 ne
rect 9975 5299 10293 5315
rect 9048 5298 9890 5299
tri 8869 5204 8963 5298 ne
tri 8963 5289 8972 5298 sw
tri 9048 5289 9057 5298 ne
rect 9057 5289 9890 5298
rect 8963 5204 8972 5289
tri 8972 5204 9057 5289 sw
tri 9057 5204 9142 5289 ne
rect 9142 5214 9890 5289
tri 9890 5214 9975 5299 sw
tri 9975 5214 10060 5299 ne
rect 10060 5279 10293 5299
tri 10293 5279 10329 5315 sw
tri 10379 5279 10415 5315 ne
rect 10415 5279 11221 5315
rect 10060 5214 10329 5279
rect 9142 5204 9975 5214
tri 8963 5110 9057 5204 ne
tri 9057 5195 9066 5204 sw
tri 9142 5195 9151 5204 ne
rect 9151 5195 9975 5204
rect 9057 5110 9066 5195
tri 9066 5110 9151 5195 sw
tri 9151 5110 9236 5195 ne
rect 9236 5154 9975 5195
tri 9975 5154 10035 5214 sw
tri 10060 5154 10120 5214 ne
rect 10120 5193 10329 5214
tri 10329 5193 10415 5279 sw
tri 10415 5193 10501 5279 ne
rect 10501 5193 11221 5279
rect 10120 5154 10415 5193
rect 9236 5110 10035 5154
tri 9057 5099 9068 5110 ne
rect 9068 5101 9151 5110
tri 9151 5101 9160 5110 sw
tri 9236 5101 9245 5110 ne
rect 9245 5101 10035 5110
rect 9068 5099 9160 5101
tri 9160 5099 9162 5101 sw
tri 9245 5099 9247 5101 ne
rect 9247 5099 10035 5101
rect 7825 5005 8645 5099
rect 7441 4979 8645 5005
tri 8645 4979 8765 5099 sw
tri 9068 5016 9151 5099 ne
rect 9151 5016 9162 5099
tri 9162 5016 9245 5099 sw
tri 9247 5016 9330 5099 ne
rect 9330 5069 10035 5099
tri 10035 5069 10120 5154 sw
tri 10120 5069 10205 5154 ne
rect 10205 5129 10415 5154
tri 10415 5129 10479 5193 sw
tri 10501 5129 10565 5193 ne
rect 10565 5129 11221 5193
rect 10205 5069 10479 5129
tri 10479 5069 10539 5129 sw
tri 10565 5069 10625 5129 ne
rect 9330 5050 10120 5069
tri 10120 5050 10139 5069 sw
tri 10205 5050 10224 5069 ne
rect 10224 5050 10539 5069
tri 10539 5050 10558 5069 sw
rect 9330 5016 10139 5050
tri 9151 4979 9188 5016 ne
rect 9188 5007 9245 5016
tri 9245 5007 9254 5016 sw
tri 9330 5007 9339 5016 ne
rect 9339 5007 10139 5016
rect 9188 4979 9254 5007
tri 4719 4846 4852 4979 ne
rect 4852 4846 5695 4979
rect 3919 4731 4131 4846
rect 3285 4690 4131 4731
rect 2757 4573 2891 4690
tri 2891 4573 3008 4690 sw
tri 3285 4573 3402 4690 ne
rect 3402 4639 4131 4690
rect 3402 4573 3683 4639
rect 2757 4503 3008 4573
rect 1864 4466 3008 4503
rect 1864 4410 2139 4466
rect 0 4333 1458 4410
rect 0 4097 294 4333
rect 530 4097 747 4333
rect 983 4097 1200 4333
rect 1436 4284 1458 4333
tri 1458 4284 1584 4410 sw
tri 1864 4284 1990 4410 ne
rect 1990 4284 2139 4410
rect 1436 4126 1584 4284
tri 1584 4126 1742 4284 sw
tri 1990 4230 2044 4284 ne
rect 2044 4230 2139 4284
rect 2375 4412 3008 4466
rect 2375 4230 2521 4412
tri 2044 4126 2148 4230 ne
rect 2148 4176 2521 4230
rect 2757 4393 3008 4412
tri 3008 4393 3188 4573 sw
tri 3402 4403 3572 4573 ne
rect 3572 4403 3683 4573
rect 3919 4610 4131 4639
rect 4367 4762 4456 4846
tri 4456 4762 4540 4846 sw
tri 4852 4762 4936 4846 ne
rect 4936 4762 5695 4846
rect 4367 4610 4540 4762
rect 3919 4573 4540 4610
tri 4540 4573 4729 4762 sw
tri 4936 4573 5125 4762 ne
rect 5125 4683 5695 4762
tri 5695 4683 5991 4979 sw
tri 6081 4683 6377 4979 ne
rect 6377 4920 7059 4979
tri 7059 4920 7118 4979 sw
tri 7441 4920 7500 4979 ne
rect 7500 4920 8765 4979
tri 8765 4920 8824 4979 sw
tri 9188 4922 9245 4979 ne
rect 9245 4922 9254 4979
tri 9254 4922 9339 5007 sw
tri 9339 4922 9424 5007 ne
rect 9424 4965 10139 5007
tri 10139 4965 10224 5050 sw
tri 10224 4965 10309 5050 ne
rect 10309 5043 10558 5050
tri 10558 5043 10565 5050 sw
rect 10309 4965 10565 5043
rect 9424 4945 10224 4965
tri 10224 4945 10244 4965 sw
tri 10309 4945 10329 4965 ne
rect 9424 4922 10244 4945
tri 9245 4920 9247 4922 ne
rect 9247 4920 9339 4922
tri 9339 4920 9341 4922 sw
tri 9424 4920 9426 4922 ne
rect 9426 4920 10244 4922
tri 10244 4920 10269 4945 sw
rect 6377 4683 7118 4920
rect 5125 4573 5991 4683
tri 5991 4573 6101 4683 sw
tri 6377 4573 6487 4683 ne
rect 6487 4673 7118 4683
tri 7118 4673 7365 4920 sw
tri 7500 4673 7747 4920 ne
rect 7747 4877 8824 4920
rect 7747 4673 7950 4877
rect 6487 4573 7365 4673
tri 7365 4573 7465 4673 sw
tri 7747 4573 7847 4673 ne
rect 7847 4641 7950 4673
rect 8186 4673 8824 4877
tri 8824 4673 9071 4920 sw
tri 9247 4828 9339 4920 ne
rect 9339 4913 9341 4920
tri 9341 4913 9348 4920 sw
tri 9426 4913 9433 4920 ne
rect 9433 4913 10269 4920
rect 9339 4828 9348 4913
tri 9348 4828 9433 4913 sw
tri 9433 4828 9518 4913 ne
rect 9518 4828 10269 4913
tri 9339 4734 9433 4828 ne
tri 9433 4819 9442 4828 sw
tri 9518 4819 9527 4828 ne
rect 9527 4819 10269 4828
rect 9433 4734 9442 4819
tri 9442 4734 9527 4819 sw
tri 9527 4734 9612 4819 ne
rect 9612 4734 10269 4819
tri 9433 4673 9494 4734 ne
rect 9494 4733 9527 4734
tri 9527 4733 9528 4734 sw
tri 9612 4733 9613 4734 ne
rect 9613 4733 10269 4734
rect 9494 4673 9528 4733
tri 9528 4673 9588 4733 sw
tri 9613 4673 9673 4733 ne
rect 8186 4641 9071 4673
rect 7847 4573 9071 4641
tri 9071 4573 9171 4673 sw
tri 9494 4640 9527 4673 ne
rect 9527 4648 9588 4673
tri 9588 4648 9613 4673 sw
rect 9527 4640 9613 4648
tri 9527 4620 9547 4640 ne
rect 3919 4519 4729 4573
rect 3919 4403 4131 4519
tri 3572 4393 3582 4403 ne
rect 3582 4393 4131 4403
rect 2757 4176 2867 4393
rect 2148 4157 2867 4176
rect 3103 4179 3188 4393
tri 3188 4179 3402 4393 sw
tri 3582 4179 3796 4393 ne
rect 3796 4283 4131 4393
rect 4367 4464 4729 4519
tri 4729 4464 4838 4573 sw
tri 5125 4497 5201 4573 ne
rect 5201 4497 6101 4573
tri 6101 4497 6177 4573 sw
tri 6487 4497 6563 4573 ne
rect 6563 4497 7465 4573
tri 7465 4497 7541 4573 sw
tri 7847 4497 7923 4573 ne
rect 7923 4497 9171 4573
tri 9171 4497 9247 4573 sw
tri 5201 4464 5234 4497 ne
rect 5234 4464 6177 4497
rect 4367 4283 4513 4464
rect 3796 4228 4513 4283
rect 4749 4228 4838 4464
rect 3796 4191 4838 4228
rect 3796 4179 4131 4191
rect 3103 4157 3402 4179
rect 2148 4126 3402 4157
rect 1436 4097 1742 4126
rect 0 4005 1742 4097
rect 0 3769 294 4005
rect 530 3769 747 4005
rect 983 3769 1200 4005
rect 1436 3769 1742 4005
rect 0 3720 1742 3769
tri 1742 3720 2148 4126 sw
tri 2148 3848 2426 4126 ne
rect 2426 4084 3402 4126
rect 2426 3848 2521 4084
rect 2757 4066 3402 4084
rect 2757 3848 2867 4066
tri 2426 3720 2554 3848 ne
rect 2554 3830 2867 3848
rect 3103 4018 3402 4066
tri 3402 4018 3563 4179 sw
tri 3796 4018 3957 4179 ne
rect 3957 4018 4131 4179
rect 3103 4011 3563 4018
rect 3103 3830 3249 4011
rect 2554 3775 3249 3830
rect 3485 3775 3563 4011
rect 2554 3738 3563 3775
rect 2554 3720 2867 3738
tri 1169 3440 1449 3720 ne
rect 1449 3440 2148 3720
tri 2148 3440 2428 3720 sw
tri 2554 3440 2834 3720 ne
rect 2834 3502 2867 3720
rect 3103 3684 3563 3738
rect 3103 3502 3249 3684
rect 2834 3448 3249 3502
rect 3485 3632 3563 3684
tri 3563 3632 3949 4018 sw
tri 3957 3955 4020 4018 ne
rect 4020 3955 4131 4018
rect 4367 4182 4838 4191
tri 4838 4182 5120 4464 sw
tri 5234 4182 5516 4464 ne
rect 5516 4297 6177 4464
tri 6177 4297 6377 4497 sw
tri 6563 4297 6763 4497 ne
rect 6763 4297 7541 4497
rect 5516 4182 6377 4297
tri 6377 4182 6492 4297 sw
tri 6763 4182 6878 4297 ne
rect 6878 4182 7541 4297
rect 4367 4137 5120 4182
rect 4367 3955 4513 4137
tri 4020 3632 4343 3955 ne
rect 4343 3901 4513 3955
rect 4749 4135 5120 4137
tri 5120 4135 5167 4182 sw
tri 5516 4135 5563 4182 ne
rect 5563 4135 6492 4182
tri 6492 4135 6539 4182 sw
tri 6878 4135 6925 4182 ne
rect 6925 4135 7541 4182
tri 7541 4135 7903 4497 sw
tri 7923 4135 8285 4497 ne
rect 8285 4455 9247 4497
rect 8285 4219 8366 4455
rect 8602 4219 8956 4455
rect 9192 4219 9247 4455
rect 8285 4135 9247 4219
rect 4749 4066 5167 4135
rect 4749 3901 4911 4066
rect 4343 3830 4911 3901
rect 5147 3830 5167 4066
rect 4343 3809 5167 3830
rect 4343 3632 4513 3809
rect 3485 3448 3628 3632
rect 2834 3440 3628 3448
rect 0 3362 1050 3440
rect 0 3126 757 3362
rect 993 3321 1050 3362
tri 1050 3321 1169 3440 sw
tri 1449 3321 1568 3440 ne
rect 1568 3383 2428 3440
tri 2428 3383 2485 3440 sw
tri 2834 3383 2891 3440 ne
rect 2891 3396 3628 3440
rect 3864 3624 3949 3632
tri 3949 3624 3957 3632 sw
tri 4343 3624 4351 3632 ne
rect 4351 3624 4513 3632
rect 3864 3440 3957 3624
tri 3957 3440 4141 3624 sw
tri 4351 3573 4402 3624 ne
rect 4402 3573 4513 3624
rect 4749 3786 5167 3809
tri 5167 3786 5516 4135 sw
tri 5563 4001 5697 4135 ne
rect 5697 4001 6539 4135
tri 6539 4001 6673 4135 sw
tri 6925 4001 7059 4135 ne
rect 7059 4115 7903 4135
tri 7903 4115 7923 4135 sw
tri 8285 4115 8305 4135 ne
rect 8305 4134 9247 4135
rect 8305 4115 8366 4134
rect 7059 4103 7923 4115
tri 7923 4103 7935 4115 sw
tri 8305 4103 8317 4115 ne
rect 7059 4001 7935 4103
tri 7935 4001 8037 4103 sw
tri 5697 3786 5912 4001 ne
rect 5912 3993 6673 4001
tri 6673 3993 6681 4001 sw
tri 7059 3993 7067 4001 ne
rect 7067 3993 8037 4001
rect 5912 3786 6681 3993
rect 4749 3739 5516 3786
rect 4749 3573 4911 3739
tri 4402 3440 4535 3573 ne
rect 4535 3503 4911 3573
rect 5147 3717 5516 3739
tri 5516 3717 5585 3786 sw
tri 5912 3717 5981 3786 ne
rect 5981 3717 6681 3786
rect 5147 3503 5585 3717
rect 4535 3440 5585 3503
rect 3864 3396 4141 3440
rect 2891 3383 4141 3396
tri 4141 3383 4198 3440 sw
tri 4535 3383 4592 3440 ne
rect 4592 3411 5585 3440
rect 4592 3383 4911 3411
rect 1568 3321 2485 3383
rect 993 3140 1169 3321
tri 1169 3140 1350 3321 sw
tri 1568 3140 1749 3321 ne
rect 1749 3246 2485 3321
tri 2485 3246 2622 3383 sw
tri 2891 3246 3028 3383 ne
rect 3028 3356 4198 3383
rect 3028 3246 3249 3356
rect 1749 3140 2622 3246
rect 993 3126 1350 3140
rect 0 2968 1350 3126
tri 1350 2968 1522 3140 sw
tri 1749 2968 1921 3140 ne
rect 1921 2977 2622 3140
tri 2622 2977 2891 3246 sw
tri 3028 3120 3154 3246 ne
rect 3154 3120 3249 3246
rect 3485 3305 4198 3356
rect 3485 3120 3628 3305
tri 3154 2977 3297 3120 ne
rect 3297 3069 3628 3120
rect 3864 3246 4198 3305
tri 4198 3246 4335 3383 sw
tri 4592 3246 4729 3383 ne
rect 4729 3246 4911 3383
rect 3864 3088 4335 3246
tri 4335 3088 4493 3246 sw
tri 4729 3088 4887 3246 ne
rect 4887 3175 4911 3246
rect 5147 3321 5585 3411
tri 5585 3321 5981 3717 sw
tri 5981 3713 5985 3717 ne
rect 5985 3713 6681 3717
tri 6681 3713 6961 3993 sw
tri 7067 3713 7347 3993 ne
rect 7347 3962 8037 3993
rect 7347 3726 7402 3962
rect 7638 3726 7750 3962
rect 7986 3726 8037 3962
tri 5985 3321 6377 3713 ne
rect 6377 3607 6961 3713
tri 6961 3607 7067 3713 sw
rect 6377 3556 7067 3607
rect 5147 3246 5981 3321
tri 5981 3246 6056 3321 sw
rect 6377 3320 6428 3556
rect 6664 3320 6782 3556
rect 7018 3320 7067 3556
rect 5147 3205 6056 3246
tri 6056 3205 6097 3246 sw
rect 5147 3175 6097 3205
rect 4887 3146 6097 3175
rect 4887 3088 5233 3146
rect 3864 3069 4493 3088
rect 3297 2977 4493 3069
rect 1921 2968 2891 2977
rect 0 2749 1151 2968
rect 0 2513 757 2749
rect 993 2732 1151 2749
rect 1387 2741 1522 2968
tri 1522 2741 1749 2968 sw
tri 1921 2808 2081 2968 ne
rect 2081 2881 2891 2968
tri 2891 2881 2987 2977 sw
tri 3297 2881 3393 2977 ne
rect 3393 2881 3628 2977
rect 2081 2808 2987 2881
tri 2987 2808 3060 2881 sw
tri 3393 2808 3466 2881 ne
rect 3466 2808 3628 2881
tri 2081 2741 2148 2808 ne
rect 2148 2741 3060 2808
tri 3060 2741 3127 2808 sw
tri 3466 2741 3533 2808 ne
rect 3533 2741 3628 2808
rect 3864 2808 4493 2977
tri 4493 2808 4773 3088 sw
tri 4887 2808 5167 3088 ne
rect 5167 2910 5233 3088
rect 5469 2910 5787 3146
rect 6023 2910 6097 3146
rect 3864 2741 4773 2808
rect 1387 2732 1749 2741
rect 993 2713 1749 2732
tri 1749 2713 1777 2741 sw
tri 2148 2713 2176 2741 ne
rect 2176 2723 3127 2741
tri 3127 2723 3145 2741 sw
tri 3533 2723 3551 2741 ne
rect 3551 2723 4773 2741
rect 2176 2713 3145 2723
rect 993 2623 1777 2713
rect 993 2513 1496 2623
rect 0 2510 1496 2513
tri 667 2230 947 2510 ne
rect 947 2387 1496 2510
rect 1732 2510 1777 2623
tri 1777 2510 1980 2713 sw
tri 2176 2510 2379 2713 ne
rect 2379 2510 3145 2713
rect 1732 2387 1980 2510
rect 947 2355 1980 2387
rect 947 2230 1151 2355
rect 0 1834 551 2230
tri 551 1834 947 2230 sw
tri 947 2119 1058 2230 ne
rect 1058 2119 1151 2230
rect 1387 2342 1980 2355
tri 1980 2342 2148 2510 sw
tri 2379 2342 2547 2510 ne
rect 2547 2342 3145 2510
rect 1387 2301 2148 2342
tri 2148 2301 2189 2342 sw
tri 2547 2301 2588 2342 ne
rect 2588 2317 3145 2342
tri 3145 2317 3551 2723 sw
tri 3551 2317 3957 2723 ne
rect 3957 2694 4773 2723
tri 4773 2694 4887 2808 sw
rect 3957 2631 4887 2694
rect 3957 2395 4011 2631
rect 4247 2395 4597 2631
rect 4833 2395 4887 2631
rect 2588 2301 3551 2317
rect 1387 2119 2189 2301
tri 1058 1834 1343 2119 ne
rect 1343 2010 2189 2119
rect 1343 1834 1496 2010
rect 0 1680 947 1834
tri 947 1680 1101 1834 sw
tri 1343 1774 1403 1834 ne
rect 1403 1774 1496 1834
rect 1732 1902 2189 2010
tri 2189 1902 2588 2301 sw
tri 2588 1902 2987 2301 ne
rect 2987 2191 3551 2301
tri 3551 2191 3677 2317 sw
rect 2987 2129 3677 2191
rect 1732 1783 2588 1902
tri 2588 1783 2707 1902 sw
rect 1732 1774 2707 1783
tri 1403 1680 1497 1774 ne
rect 1497 1721 2707 1774
rect 1497 1680 1836 1721
rect 0 1400 1101 1680
tri 1101 1400 1381 1680 sw
tri 1497 1400 1777 1680 ne
rect 1777 1485 1836 1680
rect 2072 1485 2416 1721
rect 2652 1485 2707 1721
rect 0 1284 1381 1400
tri 1381 1284 1497 1400 sw
rect 0 1225 1497 1284
rect 0 1140 470 1225
tri 0 733 407 1140 ne
rect 407 989 470 1140
rect 706 989 834 1225
rect 1070 989 1198 1225
rect 1434 989 1497 1225
rect 407 749 1497 989
rect 407 513 470 749
rect 706 513 834 749
rect 1070 513 1198 749
rect 1434 513 1497 749
rect 407 272 1497 513
rect 407 36 470 272
rect 706 36 834 272
rect 1070 36 1198 272
rect 1434 36 1497 272
rect 407 0 1497 36
rect 1777 1358 2707 1485
rect 1777 1122 1836 1358
rect 2072 1122 2416 1358
rect 2652 1122 2707 1358
rect 1777 995 2707 1122
rect 1777 759 1836 995
rect 2072 759 2416 995
rect 2652 759 2707 995
rect 1777 631 2707 759
rect 1777 395 1836 631
rect 2072 395 2416 631
rect 2652 395 2707 631
rect 1777 267 2707 395
rect 1777 31 1836 267
rect 2072 31 2416 267
rect 2652 31 2707 267
rect 1777 0 2707 31
rect 2987 1893 3037 2129
rect 3273 1893 3393 2129
rect 3629 1893 3677 2129
rect 2987 1758 3677 1893
rect 2987 1522 3037 1758
rect 3273 1522 3393 1758
rect 3629 1522 3677 1758
rect 2987 1387 3677 1522
rect 2987 1151 3037 1387
rect 3273 1151 3393 1387
rect 3629 1151 3677 1387
rect 2987 1015 3677 1151
rect 2987 779 3037 1015
rect 3273 779 3393 1015
rect 3629 779 3677 1015
rect 2987 643 3677 779
rect 2987 407 3037 643
rect 3273 407 3393 643
rect 3629 407 3677 643
rect 2987 271 3677 407
rect 2987 35 3037 271
rect 3273 35 3393 271
rect 3629 35 3677 271
rect 2987 0 3677 35
rect 3957 2295 4887 2395
rect 3957 2059 4011 2295
rect 4247 2059 4597 2295
rect 4833 2059 4887 2295
rect 3957 1959 4887 2059
rect 3957 1723 4011 1959
rect 4247 1723 4597 1959
rect 4833 1723 4887 1959
rect 3957 1623 4887 1723
rect 3957 1387 4011 1623
rect 4247 1387 4597 1623
rect 4833 1387 4887 1623
rect 3957 1287 4887 1387
rect 3957 1051 4011 1287
rect 4247 1051 4597 1287
rect 4833 1051 4887 1287
rect 3957 951 4887 1051
rect 3957 715 4011 951
rect 4247 715 4597 951
rect 4833 715 4887 951
rect 3957 615 4887 715
rect 3957 379 4011 615
rect 4247 379 4597 615
rect 4833 379 4887 615
rect 3957 279 4887 379
rect 3957 43 4011 279
rect 4247 43 4597 279
rect 4833 43 4887 279
rect 3957 0 4887 43
rect 5167 2787 6097 2910
rect 5167 2551 5233 2787
rect 5469 2551 5787 2787
rect 6023 2551 6097 2787
rect 5167 2428 6097 2551
rect 5167 2192 5233 2428
rect 5469 2192 5787 2428
rect 6023 2192 6097 2428
rect 5167 2069 6097 2192
rect 5167 1833 5233 2069
rect 5469 1833 5787 2069
rect 6023 1833 6097 2069
rect 5167 1710 6097 1833
rect 5167 1474 5233 1710
rect 5469 1474 5787 1710
rect 6023 1474 6097 1710
rect 5167 1350 6097 1474
rect 5167 1114 5233 1350
rect 5469 1114 5787 1350
rect 6023 1114 6097 1350
rect 5167 990 6097 1114
rect 5167 754 5233 990
rect 5469 754 5787 990
rect 6023 754 6097 990
rect 5167 630 6097 754
rect 5167 394 5233 630
rect 5469 394 5787 630
rect 6023 394 6097 630
rect 5167 270 6097 394
rect 5167 34 5233 270
rect 5469 34 5787 270
rect 6023 34 6097 270
rect 5167 0 6097 34
rect 6377 3228 7067 3320
rect 6377 2992 6428 3228
rect 6664 2992 6782 3228
rect 7018 2992 7067 3228
rect 6377 2900 7067 2992
rect 6377 2664 6428 2900
rect 6664 2664 6782 2900
rect 7018 2664 7067 2900
rect 6377 2572 7067 2664
rect 6377 2336 6428 2572
rect 6664 2336 6782 2572
rect 7018 2336 7067 2572
rect 6377 2244 7067 2336
rect 6377 2008 6428 2244
rect 6664 2008 6782 2244
rect 7018 2008 7067 2244
rect 6377 1916 7067 2008
rect 6377 1680 6428 1916
rect 6664 1680 6782 1916
rect 7018 1680 7067 1916
rect 6377 1588 7067 1680
rect 6377 1352 6428 1588
rect 6664 1352 6782 1588
rect 7018 1352 7067 1588
rect 6377 1260 7067 1352
rect 6377 1024 6428 1260
rect 6664 1024 6782 1260
rect 7018 1024 7067 1260
rect 6377 931 7067 1024
rect 6377 695 6428 931
rect 6664 695 6782 931
rect 7018 695 7067 931
rect 6377 602 7067 695
rect 6377 366 6428 602
rect 6664 366 6782 602
rect 7018 366 7067 602
rect 6377 273 7067 366
rect 6377 37 6428 273
rect 6664 37 6782 273
rect 7018 37 7067 273
rect 6377 0 7067 37
rect 7347 3633 8037 3726
rect 7347 3397 7402 3633
rect 7638 3397 7750 3633
rect 7986 3397 8037 3633
rect 7347 3304 8037 3397
rect 7347 3068 7402 3304
rect 7638 3068 7750 3304
rect 7986 3068 8037 3304
rect 7347 2975 8037 3068
rect 7347 2739 7402 2975
rect 7638 2739 7750 2975
rect 7986 2739 8037 2975
rect 7347 2646 8037 2739
rect 7347 2410 7402 2646
rect 7638 2410 7750 2646
rect 7986 2410 8037 2646
rect 7347 2317 8037 2410
rect 7347 2081 7402 2317
rect 7638 2081 7750 2317
rect 7986 2081 8037 2317
rect 7347 1988 8037 2081
rect 7347 1752 7402 1988
rect 7638 1752 7750 1988
rect 7986 1752 8037 1988
rect 7347 1659 8037 1752
rect 7347 1423 7402 1659
rect 7638 1423 7750 1659
rect 7986 1423 8037 1659
rect 7347 1329 8037 1423
rect 7347 1093 7402 1329
rect 7638 1093 7750 1329
rect 7986 1093 8037 1329
rect 7347 999 8037 1093
rect 7347 763 7402 999
rect 7638 763 7750 999
rect 7986 763 8037 999
rect 7347 669 8037 763
rect 7347 433 7402 669
rect 7638 433 7750 669
rect 7986 433 8037 669
rect 7347 339 8037 433
rect 7347 103 7402 339
rect 7638 103 7750 339
rect 7986 103 8037 339
rect 7347 0 8037 103
rect 8317 3898 8366 4115
rect 8602 3898 8956 4134
rect 9192 3898 9247 4134
rect 8317 3813 9247 3898
rect 8317 3577 8366 3813
rect 8602 3577 8956 3813
rect 9192 3577 9247 3813
rect 8317 3492 9247 3577
rect 8317 3256 8366 3492
rect 8602 3256 8956 3492
rect 9192 3256 9247 3492
rect 8317 3171 9247 3256
rect 8317 2935 8366 3171
rect 8602 2935 8956 3171
rect 9192 2935 9247 3171
rect 8317 2849 9247 2935
rect 8317 2613 8366 2849
rect 8602 2613 8956 2849
rect 9192 2613 9247 2849
rect 8317 2527 9247 2613
rect 8317 2291 8366 2527
rect 8602 2291 8956 2527
rect 9192 2291 9247 2527
rect 8317 2205 9247 2291
rect 8317 1969 8366 2205
rect 8602 1969 8956 2205
rect 9192 1969 9247 2205
rect 8317 1883 9247 1969
rect 8317 1647 8366 1883
rect 8602 1647 8956 1883
rect 9192 1647 9247 1883
rect 8317 1561 9247 1647
rect 8317 1325 8366 1561
rect 8602 1325 8956 1561
rect 9192 1325 9247 1561
rect 8317 1239 9247 1325
rect 8317 1003 8366 1239
rect 8602 1003 8956 1239
rect 9192 1003 9247 1239
rect 8317 917 9247 1003
rect 8317 681 8366 917
rect 8602 681 8956 917
rect 9192 681 9247 917
rect 8317 595 9247 681
rect 8317 359 8366 595
rect 8602 359 8956 595
rect 9192 359 9247 595
rect 8317 273 9247 359
rect 8317 37 8366 273
rect 8602 37 8956 273
rect 9192 37 9247 273
rect 8317 0 9247 37
rect 9547 0 9613 4640
rect 9673 0 10269 4733
rect 10329 0 10565 4965
rect 10625 0 11221 5129
rect 11281 0 11347 5368
rect 11647 5251 11703 5487
rect 11939 5251 12237 5487
rect 12473 5251 12537 5487
rect 11647 5162 12537 5251
rect 11647 4926 11703 5162
rect 11939 4926 12237 5162
rect 12473 4926 12537 5162
rect 11647 4837 12537 4926
rect 11647 4601 11703 4837
rect 11939 4601 12237 4837
rect 12473 4601 12537 4837
rect 11647 4512 12537 4601
rect 11647 4276 11703 4512
rect 11939 4276 12237 4512
rect 12473 4276 12537 4512
rect 11647 4187 12537 4276
rect 11647 3951 11703 4187
rect 11939 3951 12237 4187
rect 12473 3951 12537 4187
rect 11647 3862 12537 3951
rect 11647 3626 11703 3862
rect 11939 3626 12237 3862
rect 12473 3626 12537 3862
rect 11647 3537 12537 3626
rect 11647 3301 11703 3537
rect 11939 3301 12237 3537
rect 12473 3301 12537 3537
rect 11647 3211 12537 3301
rect 11647 2975 11703 3211
rect 11939 2975 12237 3211
rect 12473 2975 12537 3211
rect 11647 2885 12537 2975
rect 11647 2649 11703 2885
rect 11939 2649 12237 2885
rect 12473 2649 12537 2885
rect 11647 2559 12537 2649
rect 11647 2323 11703 2559
rect 11939 2323 12237 2559
rect 12473 2323 12537 2559
rect 11647 2233 12537 2323
rect 11647 1997 11703 2233
rect 11939 1997 12237 2233
rect 12473 1997 12537 2233
rect 11647 1907 12537 1997
rect 11647 1671 11703 1907
rect 11939 1671 12237 1907
rect 12473 1671 12537 1907
rect 11647 1581 12537 1671
rect 11647 1345 11703 1581
rect 11939 1345 12237 1581
rect 12473 1345 12537 1581
rect 11647 1255 12537 1345
rect 11647 1019 11703 1255
rect 11939 1019 12237 1255
rect 12473 1019 12537 1255
rect 11647 929 12537 1019
rect 11647 693 11703 929
rect 11939 693 12237 929
rect 12473 693 12537 929
rect 11647 603 12537 693
rect 11647 367 11703 603
rect 11939 367 12237 603
rect 12473 367 12537 603
rect 11647 277 12537 367
rect 11647 41 11703 277
rect 11939 41 12237 277
rect 12473 41 12537 277
rect 11647 0 12537 41
rect 12817 5948 13707 5984
rect 12817 5712 12869 5948
rect 13105 5712 13421 5948
rect 13657 5712 13707 5948
rect 12817 5617 13707 5712
rect 12817 5381 12869 5617
rect 13105 5381 13421 5617
rect 13657 5381 13707 5617
rect 12817 5286 13707 5381
rect 12817 5050 12869 5286
rect 13105 5050 13421 5286
rect 13657 5050 13707 5286
rect 12817 4955 13707 5050
rect 12817 4719 12869 4955
rect 13105 4719 13421 4955
rect 13657 4719 13707 4955
rect 12817 4624 13707 4719
rect 12817 4388 12869 4624
rect 13105 4388 13421 4624
rect 13657 4388 13707 4624
rect 12817 4293 13707 4388
rect 12817 4057 12869 4293
rect 13105 4057 13421 4293
rect 13657 4057 13707 4293
rect 12817 3962 13707 4057
rect 12817 3726 12869 3962
rect 13105 3726 13421 3962
rect 13657 3726 13707 3962
rect 12817 3631 13707 3726
rect 12817 3395 12869 3631
rect 13105 3395 13421 3631
rect 13657 3395 13707 3631
rect 12817 3300 13707 3395
rect 12817 3064 12869 3300
rect 13105 3064 13421 3300
rect 13657 3064 13707 3300
rect 12817 2969 13707 3064
rect 12817 2733 12869 2969
rect 13105 2733 13421 2969
rect 13657 2733 13707 2969
rect 12817 2638 13707 2733
rect 12817 2402 12869 2638
rect 13105 2402 13421 2638
rect 13657 2402 13707 2638
rect 12817 2307 13707 2402
rect 12817 2071 12869 2307
rect 13105 2071 13421 2307
rect 13657 2071 13707 2307
rect 12817 1976 13707 2071
rect 12817 1740 12869 1976
rect 13105 1740 13421 1976
rect 13657 1740 13707 1976
rect 12817 1644 13707 1740
rect 12817 1408 12869 1644
rect 13105 1408 13421 1644
rect 13657 1408 13707 1644
rect 12817 1312 13707 1408
rect 12817 1076 12869 1312
rect 13105 1076 13421 1312
rect 13657 1076 13707 1312
rect 12817 980 13707 1076
rect 12817 744 12869 980
rect 13105 744 13421 980
rect 13657 744 13707 980
rect 12817 648 13707 744
rect 12817 412 12869 648
rect 13105 412 13421 648
rect 13657 412 13707 648
rect 12817 316 13707 412
rect 12817 80 12869 316
rect 13105 80 13421 316
rect 13657 80 13707 316
rect 12817 0 13707 80
rect 14007 6253 14300 6489
rect 14536 6253 14624 6489
rect 14860 6253 14948 6489
rect 15184 6253 15272 6489
rect 15508 6253 15596 6489
rect 15832 6253 15920 6489
rect 16156 6253 16244 6489
rect 16480 6253 16568 6489
rect 16804 6253 16892 6489
rect 17128 6253 17216 6489
rect 17452 6253 17540 6489
rect 17776 6253 17864 6489
rect 18100 6253 18188 6489
rect 18424 6253 18512 6489
rect 18748 6253 19000 6489
rect 14007 6159 19000 6253
rect 14007 5923 14300 6159
rect 14536 5923 14624 6159
rect 14860 5923 14948 6159
rect 15184 5923 15272 6159
rect 15508 5923 15596 6159
rect 15832 5923 15920 6159
rect 16156 5923 16244 6159
rect 16480 5923 16568 6159
rect 16804 5923 16892 6159
rect 17128 5923 17216 6159
rect 17452 5923 17540 6159
rect 17776 5923 17864 6159
rect 18100 5923 18188 6159
rect 18424 5923 18512 6159
rect 18748 5923 19000 6159
rect 14007 5829 19000 5923
rect 14007 5593 14300 5829
rect 14536 5593 14624 5829
rect 14860 5593 14948 5829
rect 15184 5593 15272 5829
rect 15508 5593 15596 5829
rect 15832 5593 15920 5829
rect 16156 5593 16244 5829
rect 16480 5593 16568 5829
rect 16804 5593 16892 5829
rect 17128 5593 17216 5829
rect 17452 5593 17540 5829
rect 17776 5593 17864 5829
rect 18100 5593 18188 5829
rect 18424 5593 18512 5829
rect 18748 5593 19000 5829
rect 14007 5499 19000 5593
rect 14007 5263 14300 5499
rect 14536 5263 14624 5499
rect 14860 5263 14948 5499
rect 15184 5263 15272 5499
rect 15508 5263 15596 5499
rect 15832 5263 15920 5499
rect 16156 5263 16244 5499
rect 16480 5263 16568 5499
rect 16804 5263 16892 5499
rect 17128 5263 17216 5499
rect 17452 5263 17540 5499
rect 17776 5263 17864 5499
rect 18100 5263 18188 5499
rect 18424 5263 18512 5499
rect 18748 5263 19000 5499
rect 14007 5169 19000 5263
rect 14007 4933 14300 5169
rect 14536 4933 14624 5169
rect 14860 4933 14948 5169
rect 15184 4933 15272 5169
rect 15508 4933 15596 5169
rect 15832 4933 15920 5169
rect 16156 4933 16244 5169
rect 16480 4933 16568 5169
rect 16804 4933 16892 5169
rect 17128 4933 17216 5169
rect 17452 4933 17540 5169
rect 17776 4933 17864 5169
rect 18100 4933 18188 5169
rect 18424 4933 18512 5169
rect 18748 4933 19000 5169
rect 14007 4839 19000 4933
rect 14007 4603 14300 4839
rect 14536 4603 14624 4839
rect 14860 4603 14948 4839
rect 15184 4603 15272 4839
rect 15508 4603 15596 4839
rect 15832 4603 15920 4839
rect 16156 4603 16244 4839
rect 16480 4603 16568 4839
rect 16804 4603 16892 4839
rect 17128 4603 17216 4839
rect 17452 4603 17540 4839
rect 17776 4603 17864 4839
rect 18100 4603 18188 4839
rect 18424 4603 18512 4839
rect 18748 4603 19000 4839
rect 14007 4509 19000 4603
rect 14007 4273 14300 4509
rect 14536 4273 14624 4509
rect 14860 4273 14948 4509
rect 15184 4273 15272 4509
rect 15508 4273 15596 4509
rect 15832 4273 15920 4509
rect 16156 4273 16244 4509
rect 16480 4273 16568 4509
rect 16804 4273 16892 4509
rect 17128 4273 17216 4509
rect 17452 4273 17540 4509
rect 17776 4273 17864 4509
rect 18100 4273 18188 4509
rect 18424 4273 18512 4509
rect 18748 4273 19000 4509
rect 14007 4179 19000 4273
rect 14007 3943 14300 4179
rect 14536 3943 14624 4179
rect 14860 3943 14948 4179
rect 15184 3943 15272 4179
rect 15508 3943 15596 4179
rect 15832 3943 15920 4179
rect 16156 3943 16244 4179
rect 16480 3943 16568 4179
rect 16804 3943 16892 4179
rect 17128 3943 17216 4179
rect 17452 3943 17540 4179
rect 17776 3943 17864 4179
rect 18100 3943 18188 4179
rect 18424 3943 18512 4179
rect 18748 3943 19000 4179
rect 14007 3849 19000 3943
rect 14007 3613 14300 3849
rect 14536 3613 14624 3849
rect 14860 3613 14948 3849
rect 15184 3613 15272 3849
rect 15508 3613 15596 3849
rect 15832 3613 15920 3849
rect 16156 3613 16244 3849
rect 16480 3613 16568 3849
rect 16804 3613 16892 3849
rect 17128 3613 17216 3849
rect 17452 3613 17540 3849
rect 17776 3613 17864 3849
rect 18100 3613 18188 3849
rect 18424 3613 18512 3849
rect 18748 3613 19000 3849
rect 14007 3519 19000 3613
rect 14007 3283 14300 3519
rect 14536 3283 14624 3519
rect 14860 3283 14948 3519
rect 15184 3283 15272 3519
rect 15508 3283 15596 3519
rect 15832 3283 15920 3519
rect 16156 3283 16244 3519
rect 16480 3283 16568 3519
rect 16804 3283 16892 3519
rect 17128 3283 17216 3519
rect 17452 3283 17540 3519
rect 17776 3283 17864 3519
rect 18100 3283 18188 3519
rect 18424 3283 18512 3519
rect 18748 3283 19000 3519
rect 14007 3188 19000 3283
rect 14007 2952 14300 3188
rect 14536 2952 14624 3188
rect 14860 2952 14948 3188
rect 15184 2952 15272 3188
rect 15508 2952 15596 3188
rect 15832 2952 15920 3188
rect 16156 2952 16244 3188
rect 16480 2952 16568 3188
rect 16804 2952 16892 3188
rect 17128 2952 17216 3188
rect 17452 2952 17540 3188
rect 17776 2952 17864 3188
rect 18100 2952 18188 3188
rect 18424 2952 18512 3188
rect 18748 2952 19000 3188
rect 14007 2857 19000 2952
rect 14007 2621 14300 2857
rect 14536 2621 14624 2857
rect 14860 2621 14948 2857
rect 15184 2621 15272 2857
rect 15508 2621 15596 2857
rect 15832 2621 15920 2857
rect 16156 2621 16244 2857
rect 16480 2621 16568 2857
rect 16804 2621 16892 2857
rect 17128 2621 17216 2857
rect 17452 2621 17540 2857
rect 17776 2621 17864 2857
rect 18100 2621 18188 2857
rect 18424 2621 18512 2857
rect 18748 2621 19000 2857
rect 14007 2526 19000 2621
rect 14007 2290 14300 2526
rect 14536 2290 14624 2526
rect 14860 2290 14948 2526
rect 15184 2290 15272 2526
rect 15508 2290 15596 2526
rect 15832 2290 15920 2526
rect 16156 2290 16244 2526
rect 16480 2290 16568 2526
rect 16804 2290 16892 2526
rect 17128 2290 17216 2526
rect 17452 2290 17540 2526
rect 17776 2290 17864 2526
rect 18100 2290 18188 2526
rect 18424 2290 18512 2526
rect 18748 2290 19000 2526
rect 14007 2195 19000 2290
rect 14007 1959 14300 2195
rect 14536 1959 14624 2195
rect 14860 1959 14948 2195
rect 15184 1959 15272 2195
rect 15508 1959 15596 2195
rect 15832 1959 15920 2195
rect 16156 1959 16244 2195
rect 16480 1959 16568 2195
rect 16804 1959 16892 2195
rect 17128 1959 17216 2195
rect 17452 1959 17540 2195
rect 17776 1959 17864 2195
rect 18100 1959 18188 2195
rect 18424 1959 18512 2195
rect 18748 1959 19000 2195
rect 14007 1864 19000 1959
rect 14007 1628 14300 1864
rect 14536 1628 14624 1864
rect 14860 1628 14948 1864
rect 15184 1628 15272 1864
rect 15508 1628 15596 1864
rect 15832 1628 15920 1864
rect 16156 1628 16244 1864
rect 16480 1628 16568 1864
rect 16804 1628 16892 1864
rect 17128 1628 17216 1864
rect 17452 1628 17540 1864
rect 17776 1628 17864 1864
rect 18100 1628 18188 1864
rect 18424 1628 18512 1864
rect 18748 1628 19000 1864
rect 14007 1533 19000 1628
rect 14007 1297 14300 1533
rect 14536 1297 14624 1533
rect 14860 1297 14948 1533
rect 15184 1297 15272 1533
rect 15508 1297 15596 1533
rect 15832 1297 15920 1533
rect 16156 1297 16244 1533
rect 16480 1297 16568 1533
rect 16804 1297 16892 1533
rect 17128 1297 17216 1533
rect 17452 1297 17540 1533
rect 17776 1297 17864 1533
rect 18100 1297 18188 1533
rect 18424 1297 18512 1533
rect 18748 1297 19000 1533
rect 14007 1202 19000 1297
rect 14007 966 14300 1202
rect 14536 966 14624 1202
rect 14860 966 14948 1202
rect 15184 966 15272 1202
rect 15508 966 15596 1202
rect 15832 966 15920 1202
rect 16156 966 16244 1202
rect 16480 966 16568 1202
rect 16804 966 16892 1202
rect 17128 966 17216 1202
rect 17452 966 17540 1202
rect 17776 966 17864 1202
rect 18100 966 18188 1202
rect 18424 966 18512 1202
rect 18748 966 19000 1202
rect 14007 871 19000 966
rect 14007 635 14300 871
rect 14536 635 14624 871
rect 14860 635 14948 871
rect 15184 635 15272 871
rect 15508 635 15596 871
rect 15832 635 15920 871
rect 16156 635 16244 871
rect 16480 635 16568 871
rect 16804 635 16892 871
rect 17128 635 17216 871
rect 17452 635 17540 871
rect 17776 635 17864 871
rect 18100 635 18188 871
rect 18424 635 18512 871
rect 18748 635 19000 871
rect 14007 540 19000 635
rect 14007 304 14300 540
rect 14536 304 14624 540
rect 14860 304 14948 540
rect 15184 304 15272 540
rect 15508 304 15596 540
rect 15832 304 15920 540
rect 16156 304 16244 540
rect 16480 304 16568 540
rect 16804 304 16892 540
rect 17128 304 17216 540
rect 17452 304 17540 540
rect 17776 304 17864 540
rect 18100 304 18188 540
rect 18424 304 18512 540
rect 18748 304 19000 540
rect 14007 0 19000 304
rect 35157 8462 40000 8548
rect 35157 8226 35250 8462
rect 35486 8226 35584 8462
rect 35820 8226 35918 8462
rect 36154 8226 36252 8462
rect 36488 8226 36586 8462
rect 36822 8226 36920 8462
rect 37156 8226 37254 8462
rect 37490 8226 37588 8462
rect 37824 8226 37922 8462
rect 38158 8226 38256 8462
rect 38492 8226 38590 8462
rect 38826 8226 38924 8462
rect 39160 8226 39258 8462
rect 39494 8226 39592 8462
rect 39828 8226 40000 8462
rect 35157 8140 40000 8226
rect 35157 7904 35250 8140
rect 35486 7904 35584 8140
rect 35820 7904 35918 8140
rect 36154 7904 36252 8140
rect 36488 7904 36586 8140
rect 36822 7904 36920 8140
rect 37156 7904 37254 8140
rect 37490 7904 37588 8140
rect 37824 7904 37922 8140
rect 38158 7904 38256 8140
rect 38492 7904 38590 8140
rect 38826 7904 38924 8140
rect 39160 7904 39258 8140
rect 39494 7904 39592 8140
rect 39828 7904 40000 8140
rect 35157 7818 40000 7904
rect 35157 7582 35250 7818
rect 35486 7582 35584 7818
rect 35820 7582 35918 7818
rect 36154 7582 36252 7818
rect 36488 7582 36586 7818
rect 36822 7582 36920 7818
rect 37156 7582 37254 7818
rect 37490 7582 37588 7818
rect 37824 7582 37922 7818
rect 38158 7582 38256 7818
rect 38492 7582 38590 7818
rect 38826 7582 38924 7818
rect 39160 7582 39258 7818
rect 39494 7582 39592 7818
rect 39828 7582 40000 7818
rect 35157 7496 40000 7582
rect 35157 7260 35250 7496
rect 35486 7260 35584 7496
rect 35820 7260 35918 7496
rect 36154 7260 36252 7496
rect 36488 7260 36586 7496
rect 36822 7260 36920 7496
rect 37156 7260 37254 7496
rect 37490 7260 37588 7496
rect 37824 7260 37922 7496
rect 38158 7260 38256 7496
rect 38492 7260 38590 7496
rect 38826 7260 38924 7496
rect 39160 7260 39258 7496
rect 39494 7260 39592 7496
rect 39828 7260 40000 7496
rect 35157 7174 40000 7260
rect 35157 6938 35250 7174
rect 35486 6938 35584 7174
rect 35820 6938 35918 7174
rect 36154 6938 36252 7174
rect 36488 6938 36586 7174
rect 36822 6938 36920 7174
rect 37156 6938 37254 7174
rect 37490 6938 37588 7174
rect 37824 6938 37922 7174
rect 38158 6938 38256 7174
rect 38492 6938 38590 7174
rect 38826 6938 38924 7174
rect 39160 6938 39258 7174
rect 39494 6938 39592 7174
rect 39828 6938 40000 7174
rect 35157 6852 40000 6938
rect 35157 6616 35250 6852
rect 35486 6616 35584 6852
rect 35820 6616 35918 6852
rect 36154 6616 36252 6852
rect 36488 6616 36586 6852
rect 36822 6616 36920 6852
rect 37156 6616 37254 6852
rect 37490 6616 37588 6852
rect 37824 6616 37922 6852
rect 38158 6616 38256 6852
rect 38492 6616 38590 6852
rect 38826 6616 38924 6852
rect 39160 6616 39258 6852
rect 39494 6616 39592 6852
rect 39828 6616 40000 6852
rect 35157 6530 40000 6616
rect 35157 6294 35250 6530
rect 35486 6294 35584 6530
rect 35820 6294 35918 6530
rect 36154 6294 36252 6530
rect 36488 6294 36586 6530
rect 36822 6294 36920 6530
rect 37156 6294 37254 6530
rect 37490 6294 37588 6530
rect 37824 6294 37922 6530
rect 38158 6294 38256 6530
rect 38492 6294 38590 6530
rect 38826 6294 38924 6530
rect 39160 6294 39258 6530
rect 39494 6294 39592 6530
rect 39828 6294 40000 6530
rect 35157 6208 40000 6294
rect 35157 5972 35250 6208
rect 35486 5972 35584 6208
rect 35820 5972 35918 6208
rect 36154 5972 36252 6208
rect 36488 5972 36586 6208
rect 36822 5972 36920 6208
rect 37156 5972 37254 6208
rect 37490 5972 37588 6208
rect 37824 5972 37922 6208
rect 38158 5972 38256 6208
rect 38492 5972 38590 6208
rect 38826 5972 38924 6208
rect 39160 5972 39258 6208
rect 39494 5972 39592 6208
rect 39828 5972 40000 6208
rect 35157 5886 40000 5972
rect 35157 5650 35250 5886
rect 35486 5650 35584 5886
rect 35820 5650 35918 5886
rect 36154 5650 36252 5886
rect 36488 5650 36586 5886
rect 36822 5650 36920 5886
rect 37156 5650 37254 5886
rect 37490 5650 37588 5886
rect 37824 5650 37922 5886
rect 38158 5650 38256 5886
rect 38492 5650 38590 5886
rect 38826 5650 38924 5886
rect 39160 5650 39258 5886
rect 39494 5650 39592 5886
rect 39828 5650 40000 5886
rect 35157 5564 40000 5650
rect 35157 5328 35250 5564
rect 35486 5328 35584 5564
rect 35820 5328 35918 5564
rect 36154 5328 36252 5564
rect 36488 5328 36586 5564
rect 36822 5328 36920 5564
rect 37156 5328 37254 5564
rect 37490 5328 37588 5564
rect 37824 5328 37922 5564
rect 38158 5328 38256 5564
rect 38492 5328 38590 5564
rect 38826 5328 38924 5564
rect 39160 5328 39258 5564
rect 39494 5328 39592 5564
rect 39828 5328 40000 5564
rect 35157 5242 40000 5328
rect 35157 5006 35250 5242
rect 35486 5006 35584 5242
rect 35820 5006 35918 5242
rect 36154 5006 36252 5242
rect 36488 5006 36586 5242
rect 36822 5006 36920 5242
rect 37156 5006 37254 5242
rect 37490 5006 37588 5242
rect 37824 5006 37922 5242
rect 38158 5006 38256 5242
rect 38492 5006 38590 5242
rect 38826 5006 38924 5242
rect 39160 5006 39258 5242
rect 39494 5006 39592 5242
rect 39828 5006 40000 5242
rect 35157 4920 40000 5006
rect 35157 4684 35250 4920
rect 35486 4684 35584 4920
rect 35820 4684 35918 4920
rect 36154 4684 36252 4920
rect 36488 4684 36586 4920
rect 36822 4684 36920 4920
rect 37156 4684 37254 4920
rect 37490 4684 37588 4920
rect 37824 4684 37922 4920
rect 38158 4684 38256 4920
rect 38492 4684 38590 4920
rect 38826 4684 38924 4920
rect 39160 4684 39258 4920
rect 39494 4684 39592 4920
rect 39828 4684 40000 4920
rect 35157 4598 40000 4684
rect 35157 4362 35250 4598
rect 35486 4362 35584 4598
rect 35820 4362 35918 4598
rect 36154 4362 36252 4598
rect 36488 4362 36586 4598
rect 36822 4362 36920 4598
rect 37156 4362 37254 4598
rect 37490 4362 37588 4598
rect 37824 4362 37922 4598
rect 38158 4362 38256 4598
rect 38492 4362 38590 4598
rect 38826 4362 38924 4598
rect 39160 4362 39258 4598
rect 39494 4362 39592 4598
rect 39828 4362 40000 4598
rect 35157 4276 40000 4362
rect 35157 4040 35250 4276
rect 35486 4040 35584 4276
rect 35820 4040 35918 4276
rect 36154 4040 36252 4276
rect 36488 4040 36586 4276
rect 36822 4040 36920 4276
rect 37156 4040 37254 4276
rect 37490 4040 37588 4276
rect 37824 4040 37922 4276
rect 38158 4040 38256 4276
rect 38492 4040 38590 4276
rect 38826 4040 38924 4276
rect 39160 4040 39258 4276
rect 39494 4040 39592 4276
rect 39828 4040 40000 4276
rect 35157 3954 40000 4040
rect 35157 3718 35250 3954
rect 35486 3718 35584 3954
rect 35820 3718 35918 3954
rect 36154 3718 36252 3954
rect 36488 3718 36586 3954
rect 36822 3718 36920 3954
rect 37156 3718 37254 3954
rect 37490 3718 37588 3954
rect 37824 3718 37922 3954
rect 38158 3718 38256 3954
rect 38492 3718 38590 3954
rect 38826 3718 38924 3954
rect 39160 3718 39258 3954
rect 39494 3718 39592 3954
rect 39828 3718 40000 3954
rect 35157 3632 40000 3718
rect 35157 3396 35250 3632
rect 35486 3396 35584 3632
rect 35820 3396 35918 3632
rect 36154 3396 36252 3632
rect 36488 3396 36586 3632
rect 36822 3396 36920 3632
rect 37156 3396 37254 3632
rect 37490 3396 37588 3632
rect 37824 3396 37922 3632
rect 38158 3396 38256 3632
rect 38492 3396 38590 3632
rect 38826 3396 38924 3632
rect 39160 3396 39258 3632
rect 39494 3396 39592 3632
rect 39828 3396 40000 3632
rect 35157 3310 40000 3396
rect 35157 3074 35250 3310
rect 35486 3074 35584 3310
rect 35820 3074 35918 3310
rect 36154 3074 36252 3310
rect 36488 3074 36586 3310
rect 36822 3074 36920 3310
rect 37156 3074 37254 3310
rect 37490 3074 37588 3310
rect 37824 3074 37922 3310
rect 38158 3074 38256 3310
rect 38492 3074 38590 3310
rect 38826 3074 38924 3310
rect 39160 3074 39258 3310
rect 39494 3074 39592 3310
rect 39828 3074 40000 3310
rect 35157 2987 40000 3074
rect 35157 2751 35250 2987
rect 35486 2751 35584 2987
rect 35820 2751 35918 2987
rect 36154 2751 36252 2987
rect 36488 2751 36586 2987
rect 36822 2751 36920 2987
rect 37156 2751 37254 2987
rect 37490 2751 37588 2987
rect 37824 2751 37922 2987
rect 38158 2751 38256 2987
rect 38492 2751 38590 2987
rect 38826 2751 38924 2987
rect 39160 2751 39258 2987
rect 39494 2751 39592 2987
rect 39828 2751 40000 2987
rect 35157 2664 40000 2751
rect 35157 2428 35250 2664
rect 35486 2428 35584 2664
rect 35820 2428 35918 2664
rect 36154 2428 36252 2664
rect 36488 2428 36586 2664
rect 36822 2428 36920 2664
rect 37156 2428 37254 2664
rect 37490 2428 37588 2664
rect 37824 2428 37922 2664
rect 38158 2428 38256 2664
rect 38492 2428 38590 2664
rect 38826 2428 38924 2664
rect 39160 2428 39258 2664
rect 39494 2428 39592 2664
rect 39828 2428 40000 2664
rect 35157 2341 40000 2428
rect 35157 2105 35250 2341
rect 35486 2105 35584 2341
rect 35820 2105 35918 2341
rect 36154 2105 36252 2341
rect 36488 2105 36586 2341
rect 36822 2105 36920 2341
rect 37156 2105 37254 2341
rect 37490 2105 37588 2341
rect 37824 2105 37922 2341
rect 38158 2105 38256 2341
rect 38492 2105 38590 2341
rect 38826 2105 38924 2341
rect 39160 2105 39258 2341
rect 39494 2105 39592 2341
rect 39828 2105 40000 2341
rect 35157 2018 40000 2105
rect 35157 1782 35250 2018
rect 35486 1782 35584 2018
rect 35820 1782 35918 2018
rect 36154 1782 36252 2018
rect 36488 1782 36586 2018
rect 36822 1782 36920 2018
rect 37156 1782 37254 2018
rect 37490 1782 37588 2018
rect 37824 1782 37922 2018
rect 38158 1782 38256 2018
rect 38492 1782 38590 2018
rect 38826 1782 38924 2018
rect 39160 1782 39258 2018
rect 39494 1782 39592 2018
rect 39828 1782 40000 2018
rect 35157 1695 40000 1782
rect 35157 1459 35250 1695
rect 35486 1459 35584 1695
rect 35820 1459 35918 1695
rect 36154 1459 36252 1695
rect 36488 1459 36586 1695
rect 36822 1459 36920 1695
rect 37156 1459 37254 1695
rect 37490 1459 37588 1695
rect 37824 1459 37922 1695
rect 38158 1459 38256 1695
rect 38492 1459 38590 1695
rect 38826 1459 38924 1695
rect 39160 1459 39258 1695
rect 39494 1459 39592 1695
rect 39828 1459 40000 1695
rect 35157 1372 40000 1459
rect 35157 1136 35250 1372
rect 35486 1136 35584 1372
rect 35820 1136 35918 1372
rect 36154 1136 36252 1372
rect 36488 1136 36586 1372
rect 36822 1136 36920 1372
rect 37156 1136 37254 1372
rect 37490 1136 37588 1372
rect 37824 1136 37922 1372
rect 38158 1136 38256 1372
rect 38492 1136 38590 1372
rect 38826 1136 38924 1372
rect 39160 1136 39258 1372
rect 39494 1136 39592 1372
rect 39828 1136 40000 1372
rect 35157 1049 40000 1136
rect 35157 813 35250 1049
rect 35486 813 35584 1049
rect 35820 813 35918 1049
rect 36154 813 36252 1049
rect 36488 813 36586 1049
rect 36822 813 36920 1049
rect 37156 813 37254 1049
rect 37490 813 37588 1049
rect 37824 813 37922 1049
rect 38158 813 38256 1049
rect 38492 813 38590 1049
rect 38826 813 38924 1049
rect 39160 813 39258 1049
rect 39494 813 39592 1049
rect 39828 813 40000 1049
rect 35157 726 40000 813
rect 35157 490 35250 726
rect 35486 490 35584 726
rect 35820 490 35918 726
rect 36154 490 36252 726
rect 36488 490 36586 726
rect 36822 490 36920 726
rect 37156 490 37254 726
rect 37490 490 37588 726
rect 37824 490 37922 726
rect 38158 490 38256 726
rect 38492 490 38590 726
rect 38826 490 38924 726
rect 39160 490 39258 726
rect 39494 490 39592 726
rect 39828 490 40000 726
rect 35157 403 40000 490
rect 35157 167 35250 403
rect 35486 167 35584 403
rect 35820 167 35918 403
rect 36154 167 36252 403
rect 36488 167 36586 403
rect 36822 167 36920 403
rect 37156 167 37254 403
rect 37490 167 37588 403
rect 37824 167 37922 403
rect 38158 167 38256 403
rect 38492 167 38590 403
rect 38826 167 38924 403
rect 39160 167 39258 403
rect 39494 167 39592 403
rect 39828 167 40000 403
rect 35157 0 40000 167
<< via4 >>
rect 287 40323 523 40559
rect 610 40323 846 40559
rect 933 40323 1169 40559
rect 1256 40323 1492 40559
rect 1579 40323 1815 40559
rect 1902 40323 2138 40559
rect 2225 40323 2461 40559
rect 2548 40323 2784 40559
rect 2871 40323 3107 40559
rect 3194 40323 3430 40559
rect 3517 40323 3753 40559
rect 3840 40323 4076 40559
rect 4163 40323 4399 40559
rect 4486 40323 4722 40559
rect 4809 40323 5045 40559
rect 5132 40323 5368 40559
rect 5455 40323 5691 40559
rect 5778 40323 6014 40559
rect 6101 40323 6337 40559
rect 6424 40323 6660 40559
rect 6747 40323 6983 40559
rect 7070 40323 7306 40559
rect 7393 40323 7629 40559
rect 7716 40323 7952 40559
rect 8039 40323 8275 40559
rect 8362 40323 8598 40559
rect 8685 40323 8921 40559
rect 9008 40323 9244 40559
rect 9331 40323 9567 40559
rect 9654 40323 9890 40559
rect 9977 40323 10213 40559
rect 10300 40323 10536 40559
rect 10623 40323 10859 40559
rect 10946 40323 11182 40559
rect 11269 40323 11505 40559
rect 11592 40323 11828 40559
rect 11915 40323 12151 40559
rect 12238 40323 12474 40559
rect 12561 40323 12797 40559
rect 12884 40323 13120 40559
rect 13207 40323 13443 40559
rect 13530 40323 13766 40559
rect 13853 40323 14089 40559
rect 14176 40323 14412 40559
rect 14499 40323 14735 40559
rect 14822 40323 15058 40559
rect 15145 40323 15381 40559
rect 15468 40323 15704 40559
rect 15791 40323 16027 40559
rect 16114 40323 16350 40559
rect 16437 40323 16673 40559
rect 16760 40323 16996 40559
rect 17082 40323 17318 40559
rect 17404 40323 17640 40559
rect 17726 40323 17962 40559
rect 18048 40323 18284 40559
rect 18370 40323 18606 40559
rect 18692 40323 18928 40559
rect 19014 40323 19250 40559
rect 19336 40323 19572 40559
rect 19658 40323 19894 40559
rect 19980 40323 20216 40559
rect 20302 40323 20538 40559
rect 20624 40323 20860 40559
rect 20946 40323 21182 40559
rect 21268 40323 21504 40559
rect 21590 40323 21826 40559
rect 21912 40323 22148 40559
rect 22234 40323 22470 40559
rect 22556 40323 22792 40559
rect 22878 40323 23114 40559
rect 23200 40323 23436 40559
rect 23522 40323 23758 40559
rect 23844 40323 24080 40559
rect 24166 40323 24402 40559
rect 24488 40323 24724 40559
rect 24810 40323 25046 40559
rect 25132 40323 25368 40559
rect 287 39985 523 40221
rect 610 39985 846 40221
rect 933 39985 1169 40221
rect 1256 39985 1492 40221
rect 1579 39985 1815 40221
rect 1902 39985 2138 40221
rect 2225 39985 2461 40221
rect 2548 39985 2784 40221
rect 2871 39985 3107 40221
rect 3194 39985 3430 40221
rect 3517 39985 3753 40221
rect 3840 39985 4076 40221
rect 4163 39985 4399 40221
rect 4486 39985 4722 40221
rect 4809 39985 5045 40221
rect 5132 39985 5368 40221
rect 5455 39985 5691 40221
rect 5778 39985 6014 40221
rect 6101 39985 6337 40221
rect 6424 39985 6660 40221
rect 6747 39985 6983 40221
rect 7070 39985 7306 40221
rect 7393 39985 7629 40221
rect 7716 39985 7952 40221
rect 8039 39985 8275 40221
rect 8362 39985 8598 40221
rect 8685 39985 8921 40221
rect 9008 39985 9244 40221
rect 9331 39985 9567 40221
rect 9654 39985 9890 40221
rect 9977 39985 10213 40221
rect 10300 39985 10536 40221
rect 10623 39985 10859 40221
rect 10946 39985 11182 40221
rect 11269 39985 11505 40221
rect 11592 39985 11828 40221
rect 11915 39985 12151 40221
rect 12238 39985 12474 40221
rect 12561 39985 12797 40221
rect 12884 39985 13120 40221
rect 13207 39985 13443 40221
rect 13530 39985 13766 40221
rect 13853 39985 14089 40221
rect 14176 39985 14412 40221
rect 14499 39985 14735 40221
rect 14822 39985 15058 40221
rect 15145 39985 15381 40221
rect 15468 39985 15704 40221
rect 15791 39985 16027 40221
rect 16114 39985 16350 40221
rect 16437 39985 16673 40221
rect 16760 39985 16996 40221
rect 17082 39985 17318 40221
rect 17404 39985 17640 40221
rect 17726 39985 17962 40221
rect 18048 39985 18284 40221
rect 18370 39985 18606 40221
rect 18692 39985 18928 40221
rect 19014 39985 19250 40221
rect 19336 39985 19572 40221
rect 19658 39985 19894 40221
rect 19980 39985 20216 40221
rect 20302 39985 20538 40221
rect 20624 39985 20860 40221
rect 20946 39985 21182 40221
rect 21268 39985 21504 40221
rect 21590 39985 21826 40221
rect 21912 39985 22148 40221
rect 22234 39985 22470 40221
rect 22556 39985 22792 40221
rect 22878 39985 23114 40221
rect 23200 39985 23436 40221
rect 23522 39985 23758 40221
rect 23844 39985 24080 40221
rect 24166 39985 24402 40221
rect 24488 39985 24724 40221
rect 24810 39985 25046 40221
rect 25132 39985 25368 40221
rect 287 39647 523 39883
rect 610 39647 846 39883
rect 933 39647 1169 39883
rect 1256 39647 1492 39883
rect 1579 39647 1815 39883
rect 1902 39647 2138 39883
rect 2225 39647 2461 39883
rect 2548 39647 2784 39883
rect 2871 39647 3107 39883
rect 3194 39647 3430 39883
rect 3517 39647 3753 39883
rect 3840 39647 4076 39883
rect 4163 39647 4399 39883
rect 4486 39647 4722 39883
rect 4809 39647 5045 39883
rect 5132 39647 5368 39883
rect 5455 39647 5691 39883
rect 5778 39647 6014 39883
rect 6101 39647 6337 39883
rect 6424 39647 6660 39883
rect 6747 39647 6983 39883
rect 7070 39647 7306 39883
rect 7393 39647 7629 39883
rect 7716 39647 7952 39883
rect 8039 39647 8275 39883
rect 8362 39647 8598 39883
rect 8685 39647 8921 39883
rect 9008 39647 9244 39883
rect 9331 39647 9567 39883
rect 9654 39647 9890 39883
rect 9977 39647 10213 39883
rect 10300 39647 10536 39883
rect 10623 39647 10859 39883
rect 10946 39647 11182 39883
rect 11269 39647 11505 39883
rect 11592 39647 11828 39883
rect 11915 39647 12151 39883
rect 12238 39647 12474 39883
rect 12561 39647 12797 39883
rect 12884 39647 13120 39883
rect 13207 39647 13443 39883
rect 13530 39647 13766 39883
rect 13853 39647 14089 39883
rect 14176 39647 14412 39883
rect 14499 39647 14735 39883
rect 14822 39647 15058 39883
rect 15145 39647 15381 39883
rect 15468 39647 15704 39883
rect 15791 39647 16027 39883
rect 16114 39647 16350 39883
rect 16437 39647 16673 39883
rect 16760 39647 16996 39883
rect 17082 39647 17318 39883
rect 17404 39647 17640 39883
rect 17726 39647 17962 39883
rect 18048 39647 18284 39883
rect 18370 39647 18606 39883
rect 18692 39647 18928 39883
rect 19014 39647 19250 39883
rect 19336 39647 19572 39883
rect 19658 39647 19894 39883
rect 19980 39647 20216 39883
rect 20302 39647 20538 39883
rect 20624 39647 20860 39883
rect 20946 39647 21182 39883
rect 21268 39647 21504 39883
rect 21590 39647 21826 39883
rect 21912 39647 22148 39883
rect 22234 39647 22470 39883
rect 22556 39647 22792 39883
rect 22878 39647 23114 39883
rect 23200 39647 23436 39883
rect 23522 39647 23758 39883
rect 23844 39647 24080 39883
rect 24166 39647 24402 39883
rect 24488 39647 24724 39883
rect 24810 39647 25046 39883
rect 25132 39647 25368 39883
rect 25792 39664 26028 39900
rect 287 39309 523 39545
rect 610 39309 846 39545
rect 933 39309 1169 39545
rect 1256 39309 1492 39545
rect 1579 39309 1815 39545
rect 1902 39309 2138 39545
rect 2225 39309 2461 39545
rect 2548 39309 2784 39545
rect 2871 39309 3107 39545
rect 3194 39309 3430 39545
rect 3517 39309 3753 39545
rect 3840 39309 4076 39545
rect 4163 39309 4399 39545
rect 4486 39309 4722 39545
rect 4809 39309 5045 39545
rect 5132 39309 5368 39545
rect 5455 39309 5691 39545
rect 5778 39309 6014 39545
rect 6101 39309 6337 39545
rect 6424 39309 6660 39545
rect 6747 39309 6983 39545
rect 7070 39309 7306 39545
rect 7393 39309 7629 39545
rect 7716 39309 7952 39545
rect 8039 39309 8275 39545
rect 8362 39309 8598 39545
rect 8685 39309 8921 39545
rect 9008 39309 9244 39545
rect 9331 39309 9567 39545
rect 9654 39309 9890 39545
rect 9977 39309 10213 39545
rect 10300 39309 10536 39545
rect 10623 39309 10859 39545
rect 10946 39309 11182 39545
rect 11269 39309 11505 39545
rect 11592 39309 11828 39545
rect 11915 39309 12151 39545
rect 12238 39309 12474 39545
rect 12561 39309 12797 39545
rect 12884 39309 13120 39545
rect 13207 39309 13443 39545
rect 13530 39309 13766 39545
rect 13853 39309 14089 39545
rect 14176 39309 14412 39545
rect 14499 39309 14735 39545
rect 14822 39309 15058 39545
rect 15145 39309 15381 39545
rect 15468 39309 15704 39545
rect 15791 39309 16027 39545
rect 16114 39309 16350 39545
rect 16437 39309 16673 39545
rect 16760 39309 16996 39545
rect 17082 39309 17318 39545
rect 17404 39309 17640 39545
rect 17726 39309 17962 39545
rect 18048 39309 18284 39545
rect 18370 39309 18606 39545
rect 18692 39309 18928 39545
rect 19014 39309 19250 39545
rect 19336 39309 19572 39545
rect 19658 39309 19894 39545
rect 19980 39309 20216 39545
rect 20302 39309 20538 39545
rect 20624 39309 20860 39545
rect 20946 39309 21182 39545
rect 21268 39309 21504 39545
rect 21590 39309 21826 39545
rect 21912 39309 22148 39545
rect 22234 39309 22470 39545
rect 22556 39309 22792 39545
rect 22878 39309 23114 39545
rect 23200 39309 23436 39545
rect 23522 39309 23758 39545
rect 23844 39309 24080 39545
rect 24166 39309 24402 39545
rect 24488 39309 24724 39545
rect 24810 39309 25046 39545
rect 25132 39309 25368 39545
rect 25792 39328 26028 39564
rect 287 38971 523 39207
rect 610 38971 846 39207
rect 933 38971 1169 39207
rect 1256 38971 1492 39207
rect 1579 38971 1815 39207
rect 1902 38971 2138 39207
rect 2225 38971 2461 39207
rect 2548 38971 2784 39207
rect 2871 38971 3107 39207
rect 3194 38971 3430 39207
rect 3517 38971 3753 39207
rect 3840 38971 4076 39207
rect 4163 38971 4399 39207
rect 4486 38971 4722 39207
rect 4809 38971 5045 39207
rect 5132 38971 5368 39207
rect 5455 38971 5691 39207
rect 5778 38971 6014 39207
rect 6101 38971 6337 39207
rect 6424 38971 6660 39207
rect 6747 38971 6983 39207
rect 7070 38971 7306 39207
rect 7393 38971 7629 39207
rect 7716 38971 7952 39207
rect 8039 38971 8275 39207
rect 8362 38971 8598 39207
rect 8685 38971 8921 39207
rect 9008 38971 9244 39207
rect 9331 38971 9567 39207
rect 9654 38971 9890 39207
rect 9977 38971 10213 39207
rect 10300 38971 10536 39207
rect 10623 38971 10859 39207
rect 10946 38971 11182 39207
rect 11269 38971 11505 39207
rect 11592 38971 11828 39207
rect 11915 38971 12151 39207
rect 12238 38971 12474 39207
rect 12561 38971 12797 39207
rect 12884 38971 13120 39207
rect 13207 38971 13443 39207
rect 13530 38971 13766 39207
rect 13853 38971 14089 39207
rect 14176 38971 14412 39207
rect 14499 38971 14735 39207
rect 14822 38971 15058 39207
rect 15145 38971 15381 39207
rect 15468 38971 15704 39207
rect 15791 38971 16027 39207
rect 16114 38971 16350 39207
rect 16437 38971 16673 39207
rect 16760 38971 16996 39207
rect 17082 38971 17318 39207
rect 17404 38971 17640 39207
rect 17726 38971 17962 39207
rect 18048 38971 18284 39207
rect 18370 38971 18606 39207
rect 18692 38971 18928 39207
rect 19014 38971 19250 39207
rect 19336 38971 19572 39207
rect 19658 38971 19894 39207
rect 19980 38971 20216 39207
rect 20302 38971 20538 39207
rect 20624 38971 20860 39207
rect 20946 38971 21182 39207
rect 21268 38971 21504 39207
rect 21590 38971 21826 39207
rect 21912 38971 22148 39207
rect 22234 38971 22470 39207
rect 22556 38971 22792 39207
rect 22878 38971 23114 39207
rect 23200 38971 23436 39207
rect 23522 38971 23758 39207
rect 23844 38971 24080 39207
rect 24166 38971 24402 39207
rect 24488 38971 24724 39207
rect 24810 38971 25046 39207
rect 25132 38971 25368 39207
rect 25792 38992 26028 39228
rect 287 38633 523 38869
rect 610 38633 846 38869
rect 933 38633 1169 38869
rect 1256 38633 1492 38869
rect 1579 38633 1815 38869
rect 1902 38633 2138 38869
rect 2225 38633 2461 38869
rect 2548 38633 2784 38869
rect 2871 38633 3107 38869
rect 3194 38633 3430 38869
rect 3517 38633 3753 38869
rect 3840 38633 4076 38869
rect 4163 38633 4399 38869
rect 4486 38633 4722 38869
rect 4809 38633 5045 38869
rect 5132 38633 5368 38869
rect 5455 38633 5691 38869
rect 5778 38633 6014 38869
rect 6101 38633 6337 38869
rect 6424 38633 6660 38869
rect 6747 38633 6983 38869
rect 7070 38633 7306 38869
rect 7393 38633 7629 38869
rect 7716 38633 7952 38869
rect 8039 38633 8275 38869
rect 8362 38633 8598 38869
rect 8685 38633 8921 38869
rect 9008 38633 9244 38869
rect 9331 38633 9567 38869
rect 9654 38633 9890 38869
rect 9977 38633 10213 38869
rect 10300 38633 10536 38869
rect 10623 38633 10859 38869
rect 10946 38633 11182 38869
rect 11269 38633 11505 38869
rect 11592 38633 11828 38869
rect 11915 38633 12151 38869
rect 12238 38633 12474 38869
rect 12561 38633 12797 38869
rect 12884 38633 13120 38869
rect 13207 38633 13443 38869
rect 13530 38633 13766 38869
rect 13853 38633 14089 38869
rect 14176 38633 14412 38869
rect 14499 38633 14735 38869
rect 14822 38633 15058 38869
rect 15145 38633 15381 38869
rect 15468 38633 15704 38869
rect 15791 38633 16027 38869
rect 16114 38633 16350 38869
rect 16437 38633 16673 38869
rect 16760 38633 16996 38869
rect 17082 38633 17318 38869
rect 17404 38633 17640 38869
rect 17726 38633 17962 38869
rect 18048 38633 18284 38869
rect 18370 38633 18606 38869
rect 18692 38633 18928 38869
rect 19014 38633 19250 38869
rect 19336 38633 19572 38869
rect 19658 38633 19894 38869
rect 19980 38633 20216 38869
rect 20302 38633 20538 38869
rect 20624 38633 20860 38869
rect 20946 38633 21182 38869
rect 21268 38633 21504 38869
rect 21590 38633 21826 38869
rect 21912 38633 22148 38869
rect 22234 38633 22470 38869
rect 22556 38633 22792 38869
rect 22878 38633 23114 38869
rect 23200 38633 23436 38869
rect 23522 38633 23758 38869
rect 23844 38633 24080 38869
rect 24166 38633 24402 38869
rect 24488 38633 24724 38869
rect 24810 38633 25046 38869
rect 25132 38633 25368 38869
rect 25792 38656 26028 38892
rect 26637 38725 26873 38961
rect 287 38295 523 38531
rect 610 38295 846 38531
rect 933 38295 1169 38531
rect 1256 38295 1492 38531
rect 1579 38295 1815 38531
rect 1902 38295 2138 38531
rect 2225 38295 2461 38531
rect 2548 38295 2784 38531
rect 2871 38295 3107 38531
rect 3194 38295 3430 38531
rect 3517 38295 3753 38531
rect 3840 38295 4076 38531
rect 4163 38295 4399 38531
rect 4486 38295 4722 38531
rect 4809 38295 5045 38531
rect 5132 38295 5368 38531
rect 5455 38295 5691 38531
rect 5778 38295 6014 38531
rect 6101 38295 6337 38531
rect 6424 38295 6660 38531
rect 6747 38295 6983 38531
rect 7070 38295 7306 38531
rect 7393 38295 7629 38531
rect 7716 38295 7952 38531
rect 8039 38295 8275 38531
rect 8362 38295 8598 38531
rect 8685 38295 8921 38531
rect 9008 38295 9244 38531
rect 9331 38295 9567 38531
rect 9654 38295 9890 38531
rect 9977 38295 10213 38531
rect 10300 38295 10536 38531
rect 10623 38295 10859 38531
rect 10946 38295 11182 38531
rect 11269 38295 11505 38531
rect 11592 38295 11828 38531
rect 11915 38295 12151 38531
rect 12238 38295 12474 38531
rect 12561 38295 12797 38531
rect 12884 38295 13120 38531
rect 13207 38295 13443 38531
rect 13530 38295 13766 38531
rect 13853 38295 14089 38531
rect 14176 38295 14412 38531
rect 14499 38295 14735 38531
rect 14822 38295 15058 38531
rect 15145 38295 15381 38531
rect 15468 38295 15704 38531
rect 15791 38295 16027 38531
rect 16114 38295 16350 38531
rect 16437 38295 16673 38531
rect 16760 38295 16996 38531
rect 17082 38295 17318 38531
rect 17404 38295 17640 38531
rect 17726 38295 17962 38531
rect 18048 38295 18284 38531
rect 18370 38295 18606 38531
rect 18692 38295 18928 38531
rect 19014 38295 19250 38531
rect 19336 38295 19572 38531
rect 19658 38295 19894 38531
rect 19980 38295 20216 38531
rect 20302 38295 20538 38531
rect 20624 38295 20860 38531
rect 20946 38295 21182 38531
rect 21268 38295 21504 38531
rect 21590 38295 21826 38531
rect 21912 38295 22148 38531
rect 22234 38295 22470 38531
rect 22556 38295 22792 38531
rect 22878 38295 23114 38531
rect 23200 38295 23436 38531
rect 23522 38295 23758 38531
rect 23844 38295 24080 38531
rect 24166 38295 24402 38531
rect 24488 38295 24724 38531
rect 24810 38295 25046 38531
rect 25132 38295 25368 38531
rect 25792 38320 26028 38556
rect 26637 38389 26873 38625
rect 287 37957 523 38193
rect 610 37957 846 38193
rect 933 37957 1169 38193
rect 1256 37957 1492 38193
rect 1579 37957 1815 38193
rect 1902 37957 2138 38193
rect 2225 37957 2461 38193
rect 2548 37957 2784 38193
rect 2871 37957 3107 38193
rect 3194 37957 3430 38193
rect 3517 37957 3753 38193
rect 3840 37957 4076 38193
rect 4163 37957 4399 38193
rect 4486 37957 4722 38193
rect 4809 37957 5045 38193
rect 5132 37957 5368 38193
rect 5455 37957 5691 38193
rect 5778 37957 6014 38193
rect 6101 37957 6337 38193
rect 6424 37957 6660 38193
rect 6747 37957 6983 38193
rect 7070 37957 7306 38193
rect 7393 37957 7629 38193
rect 7716 37957 7952 38193
rect 8039 37957 8275 38193
rect 8362 37957 8598 38193
rect 8685 37957 8921 38193
rect 9008 37957 9244 38193
rect 9331 37957 9567 38193
rect 9654 37957 9890 38193
rect 9977 37957 10213 38193
rect 10300 37957 10536 38193
rect 10623 37957 10859 38193
rect 10946 37957 11182 38193
rect 11269 37957 11505 38193
rect 11592 37957 11828 38193
rect 11915 37957 12151 38193
rect 12238 37957 12474 38193
rect 12561 37957 12797 38193
rect 12884 37957 13120 38193
rect 13207 37957 13443 38193
rect 13530 37957 13766 38193
rect 13853 37957 14089 38193
rect 14176 37957 14412 38193
rect 14499 37957 14735 38193
rect 14822 37957 15058 38193
rect 15145 37957 15381 38193
rect 15468 37957 15704 38193
rect 15791 37957 16027 38193
rect 16114 37957 16350 38193
rect 16437 37957 16673 38193
rect 16760 37957 16996 38193
rect 17082 37957 17318 38193
rect 17404 37957 17640 38193
rect 17726 37957 17962 38193
rect 18048 37957 18284 38193
rect 18370 37957 18606 38193
rect 18692 37957 18928 38193
rect 19014 37957 19250 38193
rect 19336 37957 19572 38193
rect 19658 37957 19894 38193
rect 19980 37957 20216 38193
rect 20302 37957 20538 38193
rect 20624 37957 20860 38193
rect 20946 37957 21182 38193
rect 21268 37957 21504 38193
rect 21590 37957 21826 38193
rect 21912 37957 22148 38193
rect 22234 37957 22470 38193
rect 22556 37957 22792 38193
rect 22878 37957 23114 38193
rect 23200 37957 23436 38193
rect 23522 37957 23758 38193
rect 23844 37957 24080 38193
rect 24166 37957 24402 38193
rect 24488 37957 24724 38193
rect 24810 37957 25046 38193
rect 25132 37957 25368 38193
rect 25792 37984 26028 38220
rect 26637 38053 26873 38289
rect 27393 38063 27629 38299
rect 287 37619 523 37855
rect 610 37619 846 37855
rect 933 37619 1169 37855
rect 1256 37619 1492 37855
rect 1579 37619 1815 37855
rect 1902 37619 2138 37855
rect 2225 37619 2461 37855
rect 2548 37619 2784 37855
rect 2871 37619 3107 37855
rect 3194 37619 3430 37855
rect 3517 37619 3753 37855
rect 3840 37619 4076 37855
rect 4163 37619 4399 37855
rect 4486 37619 4722 37855
rect 4809 37619 5045 37855
rect 5132 37619 5368 37855
rect 5455 37619 5691 37855
rect 5778 37619 6014 37855
rect 6101 37619 6337 37855
rect 6424 37619 6660 37855
rect 6747 37619 6983 37855
rect 7070 37619 7306 37855
rect 7393 37619 7629 37855
rect 7716 37619 7952 37855
rect 8039 37619 8275 37855
rect 8362 37619 8598 37855
rect 8685 37619 8921 37855
rect 9008 37619 9244 37855
rect 9331 37619 9567 37855
rect 9654 37619 9890 37855
rect 9977 37619 10213 37855
rect 10300 37619 10536 37855
rect 10623 37619 10859 37855
rect 10946 37619 11182 37855
rect 11269 37619 11505 37855
rect 11592 37619 11828 37855
rect 11915 37619 12151 37855
rect 12238 37619 12474 37855
rect 12561 37619 12797 37855
rect 12884 37619 13120 37855
rect 13207 37619 13443 37855
rect 13530 37619 13766 37855
rect 13853 37619 14089 37855
rect 14176 37619 14412 37855
rect 14499 37619 14735 37855
rect 14822 37619 15058 37855
rect 15145 37619 15381 37855
rect 15468 37619 15704 37855
rect 15791 37619 16027 37855
rect 16114 37619 16350 37855
rect 16437 37619 16673 37855
rect 16760 37619 16996 37855
rect 17082 37619 17318 37855
rect 17404 37619 17640 37855
rect 17726 37619 17962 37855
rect 18048 37619 18284 37855
rect 18370 37619 18606 37855
rect 18692 37619 18928 37855
rect 19014 37619 19250 37855
rect 19336 37619 19572 37855
rect 19658 37619 19894 37855
rect 19980 37619 20216 37855
rect 20302 37619 20538 37855
rect 20624 37619 20860 37855
rect 20946 37619 21182 37855
rect 21268 37619 21504 37855
rect 21590 37619 21826 37855
rect 21912 37619 22148 37855
rect 22234 37619 22470 37855
rect 22556 37619 22792 37855
rect 22878 37619 23114 37855
rect 23200 37619 23436 37855
rect 23522 37619 23758 37855
rect 23844 37619 24080 37855
rect 24166 37619 24402 37855
rect 24488 37619 24724 37855
rect 24810 37619 25046 37855
rect 25132 37619 25368 37855
rect 25792 37648 26028 37884
rect 26637 37717 26873 37953
rect 27393 37727 27629 37963
rect 287 37281 523 37517
rect 610 37281 846 37517
rect 933 37281 1169 37517
rect 1256 37281 1492 37517
rect 1579 37281 1815 37517
rect 1902 37281 2138 37517
rect 2225 37281 2461 37517
rect 2548 37281 2784 37517
rect 2871 37281 3107 37517
rect 3194 37281 3430 37517
rect 3517 37281 3753 37517
rect 3840 37281 4076 37517
rect 4163 37281 4399 37517
rect 4486 37281 4722 37517
rect 4809 37281 5045 37517
rect 5132 37281 5368 37517
rect 5455 37281 5691 37517
rect 5778 37281 6014 37517
rect 6101 37281 6337 37517
rect 6424 37281 6660 37517
rect 6747 37281 6983 37517
rect 7070 37281 7306 37517
rect 7393 37281 7629 37517
rect 7716 37281 7952 37517
rect 8039 37281 8275 37517
rect 8362 37281 8598 37517
rect 8685 37281 8921 37517
rect 9008 37281 9244 37517
rect 9331 37281 9567 37517
rect 9654 37281 9890 37517
rect 9977 37281 10213 37517
rect 10300 37281 10536 37517
rect 10623 37281 10859 37517
rect 10946 37281 11182 37517
rect 11269 37281 11505 37517
rect 11592 37281 11828 37517
rect 11915 37281 12151 37517
rect 12238 37281 12474 37517
rect 12561 37281 12797 37517
rect 12884 37281 13120 37517
rect 13207 37281 13443 37517
rect 13530 37281 13766 37517
rect 13853 37281 14089 37517
rect 14176 37281 14412 37517
rect 14499 37281 14735 37517
rect 14822 37281 15058 37517
rect 15145 37281 15381 37517
rect 15468 37281 15704 37517
rect 15791 37281 16027 37517
rect 16114 37281 16350 37517
rect 16437 37281 16673 37517
rect 16760 37281 16996 37517
rect 17082 37281 17318 37517
rect 17404 37281 17640 37517
rect 17726 37281 17962 37517
rect 18048 37281 18284 37517
rect 18370 37281 18606 37517
rect 18692 37281 18928 37517
rect 19014 37281 19250 37517
rect 19336 37281 19572 37517
rect 19658 37281 19894 37517
rect 19980 37281 20216 37517
rect 20302 37281 20538 37517
rect 20624 37281 20860 37517
rect 20946 37281 21182 37517
rect 21268 37281 21504 37517
rect 21590 37281 21826 37517
rect 21912 37281 22148 37517
rect 22234 37281 22470 37517
rect 22556 37281 22792 37517
rect 22878 37281 23114 37517
rect 23200 37281 23436 37517
rect 23522 37281 23758 37517
rect 23844 37281 24080 37517
rect 24166 37281 24402 37517
rect 24488 37281 24724 37517
rect 24810 37281 25046 37517
rect 25132 37281 25368 37517
rect 25792 37312 26028 37548
rect 26637 37381 26873 37617
rect 27393 37391 27629 37627
rect 287 36943 523 37179
rect 610 36943 846 37179
rect 933 36943 1169 37179
rect 1256 36943 1492 37179
rect 1579 36943 1815 37179
rect 1902 36943 2138 37179
rect 2225 36943 2461 37179
rect 2548 36943 2784 37179
rect 2871 36943 3107 37179
rect 3194 36943 3430 37179
rect 3517 36943 3753 37179
rect 3840 36943 4076 37179
rect 4163 36943 4399 37179
rect 4486 36943 4722 37179
rect 4809 36943 5045 37179
rect 5132 36943 5368 37179
rect 5455 36943 5691 37179
rect 5778 36943 6014 37179
rect 6101 36943 6337 37179
rect 6424 36943 6660 37179
rect 6747 36943 6983 37179
rect 7070 36943 7306 37179
rect 7393 36943 7629 37179
rect 7716 36943 7952 37179
rect 8039 36943 8275 37179
rect 8362 36943 8598 37179
rect 8685 36943 8921 37179
rect 9008 36943 9244 37179
rect 9331 36943 9567 37179
rect 9654 36943 9890 37179
rect 9977 36943 10213 37179
rect 10300 36943 10536 37179
rect 10623 36943 10859 37179
rect 10946 36943 11182 37179
rect 11269 36943 11505 37179
rect 11592 36943 11828 37179
rect 11915 36943 12151 37179
rect 12238 36943 12474 37179
rect 12561 36943 12797 37179
rect 12884 36943 13120 37179
rect 13207 36943 13443 37179
rect 13530 36943 13766 37179
rect 13853 36943 14089 37179
rect 14176 36943 14412 37179
rect 14499 36943 14735 37179
rect 14822 36943 15058 37179
rect 15145 36943 15381 37179
rect 15468 36943 15704 37179
rect 15791 36943 16027 37179
rect 16114 36943 16350 37179
rect 16437 36943 16673 37179
rect 16760 36943 16996 37179
rect 17082 36943 17318 37179
rect 17404 36943 17640 37179
rect 17726 36943 17962 37179
rect 18048 36943 18284 37179
rect 18370 36943 18606 37179
rect 18692 36943 18928 37179
rect 19014 36943 19250 37179
rect 19336 36943 19572 37179
rect 19658 36943 19894 37179
rect 19980 36943 20216 37179
rect 20302 36943 20538 37179
rect 20624 36943 20860 37179
rect 20946 36943 21182 37179
rect 21268 36943 21504 37179
rect 21590 36943 21826 37179
rect 21912 36943 22148 37179
rect 22234 36943 22470 37179
rect 22556 36943 22792 37179
rect 22878 36943 23114 37179
rect 23200 36943 23436 37179
rect 23522 36943 23758 37179
rect 23844 36943 24080 37179
rect 24166 36943 24402 37179
rect 24488 36943 24724 37179
rect 24810 36943 25046 37179
rect 25132 36943 25368 37179
rect 25792 36975 26028 37211
rect 26637 37045 26873 37281
rect 27393 37055 27629 37291
rect 28238 37124 28474 37360
rect 287 36605 523 36841
rect 610 36605 846 36841
rect 933 36605 1169 36841
rect 1256 36605 1492 36841
rect 1579 36605 1815 36841
rect 1902 36605 2138 36841
rect 2225 36605 2461 36841
rect 2548 36605 2784 36841
rect 2871 36605 3107 36841
rect 3194 36605 3430 36841
rect 3517 36605 3753 36841
rect 3840 36605 4076 36841
rect 4163 36605 4399 36841
rect 4486 36605 4722 36841
rect 4809 36605 5045 36841
rect 5132 36605 5368 36841
rect 5455 36605 5691 36841
rect 5778 36605 6014 36841
rect 6101 36605 6337 36841
rect 6424 36605 6660 36841
rect 6747 36605 6983 36841
rect 7070 36605 7306 36841
rect 7393 36605 7629 36841
rect 7716 36605 7952 36841
rect 8039 36605 8275 36841
rect 8362 36605 8598 36841
rect 8685 36605 8921 36841
rect 9008 36605 9244 36841
rect 9331 36605 9567 36841
rect 9654 36605 9890 36841
rect 9977 36605 10213 36841
rect 10300 36605 10536 36841
rect 10623 36605 10859 36841
rect 10946 36605 11182 36841
rect 11269 36605 11505 36841
rect 11592 36605 11828 36841
rect 11915 36605 12151 36841
rect 12238 36605 12474 36841
rect 12561 36605 12797 36841
rect 12884 36605 13120 36841
rect 13207 36605 13443 36841
rect 13530 36605 13766 36841
rect 13853 36605 14089 36841
rect 14176 36605 14412 36841
rect 14499 36605 14735 36841
rect 14822 36605 15058 36841
rect 15145 36605 15381 36841
rect 15468 36605 15704 36841
rect 15791 36605 16027 36841
rect 16114 36605 16350 36841
rect 16437 36605 16673 36841
rect 16760 36605 16996 36841
rect 17082 36605 17318 36841
rect 17404 36605 17640 36841
rect 17726 36605 17962 36841
rect 18048 36605 18284 36841
rect 18370 36605 18606 36841
rect 18692 36605 18928 36841
rect 19014 36605 19250 36841
rect 19336 36605 19572 36841
rect 19658 36605 19894 36841
rect 19980 36605 20216 36841
rect 20302 36605 20538 36841
rect 20624 36605 20860 36841
rect 20946 36605 21182 36841
rect 21268 36605 21504 36841
rect 21590 36605 21826 36841
rect 21912 36605 22148 36841
rect 22234 36605 22470 36841
rect 22556 36605 22792 36841
rect 22878 36605 23114 36841
rect 23200 36605 23436 36841
rect 23522 36605 23758 36841
rect 23844 36605 24080 36841
rect 24166 36605 24402 36841
rect 24488 36605 24724 36841
rect 24810 36605 25046 36841
rect 25132 36605 25368 36841
rect 25792 36638 26028 36874
rect 26637 36709 26873 36945
rect 27393 36719 27629 36955
rect 28238 36788 28474 37024
rect 287 36267 523 36503
rect 610 36267 846 36503
rect 933 36267 1169 36503
rect 1256 36267 1492 36503
rect 1579 36267 1815 36503
rect 1902 36267 2138 36503
rect 2225 36267 2461 36503
rect 2548 36267 2784 36503
rect 2871 36267 3107 36503
rect 3194 36267 3430 36503
rect 3517 36267 3753 36503
rect 3840 36267 4076 36503
rect 4163 36267 4399 36503
rect 4486 36267 4722 36503
rect 4809 36267 5045 36503
rect 5132 36267 5368 36503
rect 5455 36267 5691 36503
rect 5778 36267 6014 36503
rect 6101 36267 6337 36503
rect 6424 36267 6660 36503
rect 6747 36267 6983 36503
rect 7070 36267 7306 36503
rect 7393 36267 7629 36503
rect 7716 36267 7952 36503
rect 8039 36267 8275 36503
rect 8362 36267 8598 36503
rect 8685 36267 8921 36503
rect 9008 36267 9244 36503
rect 9331 36267 9567 36503
rect 9654 36267 9890 36503
rect 9977 36267 10213 36503
rect 10300 36267 10536 36503
rect 10623 36267 10859 36503
rect 10946 36267 11182 36503
rect 11269 36267 11505 36503
rect 11592 36267 11828 36503
rect 11915 36267 12151 36503
rect 12238 36267 12474 36503
rect 12561 36267 12797 36503
rect 12884 36267 13120 36503
rect 13207 36267 13443 36503
rect 13530 36267 13766 36503
rect 13853 36267 14089 36503
rect 14176 36267 14412 36503
rect 14499 36267 14735 36503
rect 14822 36267 15058 36503
rect 15145 36267 15381 36503
rect 15468 36267 15704 36503
rect 15791 36267 16027 36503
rect 16114 36267 16350 36503
rect 16437 36267 16673 36503
rect 16760 36267 16996 36503
rect 17082 36267 17318 36503
rect 17404 36267 17640 36503
rect 17726 36267 17962 36503
rect 18048 36267 18284 36503
rect 18370 36267 18606 36503
rect 18692 36267 18928 36503
rect 19014 36267 19250 36503
rect 19336 36267 19572 36503
rect 19658 36267 19894 36503
rect 19980 36267 20216 36503
rect 20302 36267 20538 36503
rect 20624 36267 20860 36503
rect 20946 36267 21182 36503
rect 21268 36267 21504 36503
rect 21590 36267 21826 36503
rect 21912 36267 22148 36503
rect 22234 36267 22470 36503
rect 22556 36267 22792 36503
rect 22878 36267 23114 36503
rect 23200 36267 23436 36503
rect 23522 36267 23758 36503
rect 23844 36267 24080 36503
rect 24166 36267 24402 36503
rect 24488 36267 24724 36503
rect 24810 36267 25046 36503
rect 25132 36267 25368 36503
rect 25792 36301 26028 36537
rect 26637 36373 26873 36609
rect 27393 36383 27629 36619
rect 28238 36452 28474 36688
rect 28994 36462 29230 36698
rect 287 35929 523 36165
rect 610 35929 846 36165
rect 933 35929 1169 36165
rect 1256 35929 1492 36165
rect 1579 35929 1815 36165
rect 1902 35929 2138 36165
rect 2225 35929 2461 36165
rect 2548 35929 2784 36165
rect 2871 35929 3107 36165
rect 3194 35929 3430 36165
rect 3517 35929 3753 36165
rect 3840 35929 4076 36165
rect 4163 35929 4399 36165
rect 4486 35929 4722 36165
rect 4809 35929 5045 36165
rect 5132 35929 5368 36165
rect 5455 35929 5691 36165
rect 5778 35929 6014 36165
rect 6101 35929 6337 36165
rect 6424 35929 6660 36165
rect 6747 35929 6983 36165
rect 7070 35929 7306 36165
rect 7393 35929 7629 36165
rect 7716 35929 7952 36165
rect 8039 35929 8275 36165
rect 8362 35929 8598 36165
rect 8685 35929 8921 36165
rect 9008 35929 9244 36165
rect 9331 35929 9567 36165
rect 9654 35929 9890 36165
rect 9977 35929 10213 36165
rect 10300 35929 10536 36165
rect 10623 35929 10859 36165
rect 10946 35929 11182 36165
rect 11269 35929 11505 36165
rect 11592 35929 11828 36165
rect 11915 35929 12151 36165
rect 12238 35929 12474 36165
rect 12561 35929 12797 36165
rect 12884 35929 13120 36165
rect 13207 35929 13443 36165
rect 13530 35929 13766 36165
rect 13853 35929 14089 36165
rect 14176 35929 14412 36165
rect 14499 35929 14735 36165
rect 14822 35929 15058 36165
rect 15145 35929 15381 36165
rect 15468 35929 15704 36165
rect 15791 35929 16027 36165
rect 16114 35929 16350 36165
rect 16437 35929 16673 36165
rect 16760 35929 16996 36165
rect 17082 35929 17318 36165
rect 17404 35929 17640 36165
rect 17726 35929 17962 36165
rect 18048 35929 18284 36165
rect 18370 35929 18606 36165
rect 18692 35929 18928 36165
rect 19014 35929 19250 36165
rect 19336 35929 19572 36165
rect 19658 35929 19894 36165
rect 19980 35929 20216 36165
rect 20302 35929 20538 36165
rect 20624 35929 20860 36165
rect 20946 35929 21182 36165
rect 21268 35929 21504 36165
rect 21590 35929 21826 36165
rect 21912 35929 22148 36165
rect 22234 35929 22470 36165
rect 22556 35929 22792 36165
rect 22878 35929 23114 36165
rect 23200 35929 23436 36165
rect 23522 35929 23758 36165
rect 23844 35929 24080 36165
rect 24166 35929 24402 36165
rect 24488 35929 24724 36165
rect 24810 35929 25046 36165
rect 25132 35929 25368 36165
rect 25792 35964 26028 36200
rect 26637 36036 26873 36272
rect 27393 36047 27629 36283
rect 28238 36116 28474 36352
rect 28994 36126 29230 36362
rect 25792 35627 26028 35863
rect 26637 35699 26873 35935
rect 27393 35711 27629 35947
rect 28238 35780 28474 36016
rect 28994 35790 29230 36026
rect 25792 35290 26028 35526
rect 26637 35362 26873 35598
rect 27393 35374 27629 35610
rect 28238 35444 28474 35680
rect 28994 35454 29230 35690
rect 29839 35523 30075 35759
rect 25792 34953 26028 35189
rect 26637 35025 26873 35261
rect 27393 35037 27629 35273
rect 28238 35108 28474 35344
rect 28994 35118 29230 35354
rect 29839 35187 30075 35423
rect 25792 34616 26028 34852
rect 26637 34688 26873 34924
rect 27393 34700 27629 34936
rect 28238 34772 28474 35008
rect 28994 34782 29230 35018
rect 29839 34851 30075 35087
rect 30595 34861 30831 35097
rect 25792 34279 26028 34515
rect 26637 34351 26873 34587
rect 27393 34363 27629 34599
rect 28238 34435 28474 34671
rect 28994 34446 29230 34682
rect 29839 34515 30075 34751
rect 30595 34525 30831 34761
rect 25792 33942 26028 34178
rect 26637 34014 26873 34250
rect 27393 34026 27629 34262
rect 28238 34098 28474 34334
rect 28994 34110 29230 34346
rect 29839 34179 30075 34415
rect 30595 34189 30831 34425
rect 25792 33605 26028 33841
rect 26637 33677 26873 33913
rect 27393 33689 27629 33925
rect 28238 33761 28474 33997
rect 28994 33773 29230 34009
rect 29839 33843 30075 34079
rect 30595 33853 30831 34089
rect 31440 33922 31676 34158
rect 26637 33340 26873 33576
rect 27393 33352 27629 33588
rect 28238 33424 28474 33660
rect 28994 33436 29230 33672
rect 29839 33507 30075 33743
rect 30595 33517 30831 33753
rect 31440 33586 31676 33822
rect 26637 33003 26873 33239
rect 27393 33015 27629 33251
rect 28238 33087 28474 33323
rect 28994 33099 29230 33335
rect 29839 33171 30075 33407
rect 30595 33181 30831 33417
rect 31440 33250 31676 33486
rect 32119 33337 32355 33573
rect 26637 32666 26873 32902
rect 27393 32678 27629 32914
rect 28238 32750 28474 32986
rect 28994 32762 29230 32998
rect 29839 32834 30075 33070
rect 30595 32845 30831 33081
rect 31440 32914 31676 33150
rect 32119 33001 32355 33237
rect 27393 32341 27629 32577
rect 28238 32413 28474 32649
rect 28994 32425 29230 32661
rect 29839 32497 30075 32733
rect 30595 32509 30831 32745
rect 31440 32578 31676 32814
rect 32119 32665 32355 32901
rect 27393 32004 27629 32240
rect 28238 32076 28474 32312
rect 28994 32088 29230 32324
rect 29839 32160 30075 32396
rect 30595 32172 30831 32408
rect 31440 32242 31676 32478
rect 32119 32329 32355 32565
rect 32964 32398 33200 32634
rect 28238 31739 28474 31975
rect 28994 31751 29230 31987
rect 29839 31823 30075 32059
rect 30595 31835 30831 32071
rect 31440 31906 31676 32142
rect 32119 31993 32355 32229
rect 32964 32062 33200 32298
rect 28238 31402 28474 31638
rect 28994 31414 29230 31650
rect 29839 31486 30075 31722
rect 30595 31498 30831 31734
rect 31440 31570 31676 31806
rect 32119 31657 32355 31893
rect 32964 31726 33200 31962
rect 33720 31736 33956 31972
rect 28238 31065 28474 31301
rect 28994 31077 29230 31313
rect 29839 31149 30075 31385
rect 30595 31161 30831 31397
rect 31440 31233 31676 31469
rect 32119 31321 32355 31557
rect 32964 31390 33200 31626
rect 33720 31400 33956 31636
rect 28994 30740 29230 30976
rect 29839 30812 30075 31048
rect 30595 30824 30831 31060
rect 31440 30896 31676 31132
rect 32119 30985 32355 31221
rect 32964 31054 33200 31290
rect 33720 31064 33956 31300
rect 28994 30403 29230 30639
rect 29839 30475 30075 30711
rect 30595 30487 30831 30723
rect 31440 30559 31676 30795
rect 32119 30648 32355 30884
rect 32964 30718 33200 30954
rect 33720 30728 33956 30964
rect 34565 30797 34801 31033
rect 29839 30138 30075 30374
rect 30595 30150 30831 30386
rect 31440 30222 31676 30458
rect 32119 30311 32355 30547
rect 32964 30382 33200 30618
rect 33720 30392 33956 30628
rect 34565 30461 34801 30697
rect 29839 29801 30075 30037
rect 30595 29813 30831 30049
rect 31440 29885 31676 30121
rect 32119 29974 32355 30210
rect 32964 30046 33200 30282
rect 33720 30056 33956 30292
rect 34565 30125 34801 30361
rect 29839 29464 30075 29700
rect 30595 29476 30831 29712
rect 31440 29548 31676 29784
rect 32119 29637 32355 29873
rect 32964 29709 33200 29945
rect 33720 29720 33956 29956
rect 34565 29789 34801 30025
rect 35365 29997 35601 30233
rect 30595 29139 30831 29375
rect 31440 29211 31676 29447
rect 32119 29300 32355 29536
rect 32964 29372 33200 29608
rect 33720 29384 33956 29620
rect 34565 29453 34801 29689
rect 35365 29665 35601 29901
rect 30595 28802 30831 29038
rect 31440 28874 31676 29110
rect 32119 28963 32355 29199
rect 32964 29035 33200 29271
rect 33720 29047 33956 29283
rect 34565 29117 34801 29353
rect 35365 29333 35601 29569
rect 31440 28537 31676 28773
rect 32119 28626 32355 28862
rect 32964 28698 33200 28934
rect 33720 28710 33956 28946
rect 34565 28781 34801 29017
rect 35365 29001 35601 29237
rect 36237 29125 36473 29361
rect 31440 28200 31676 28436
rect 32119 28289 32355 28525
rect 32964 28361 33200 28597
rect 33720 28373 33956 28609
rect 34565 28445 34801 28681
rect 35365 28669 35601 28905
rect 36237 28793 36473 29029
rect 31440 27863 31676 28099
rect 32119 27952 32355 28188
rect 32964 28024 33200 28260
rect 33720 28036 33956 28272
rect 34565 28108 34801 28344
rect 35365 28337 35601 28573
rect 36237 28461 36473 28697
rect 32119 27615 32355 27851
rect 32964 27687 33200 27923
rect 33720 27699 33956 27935
rect 34565 27771 34801 28007
rect 35365 28005 35601 28241
rect 36237 28129 36473 28365
rect 37123 28239 37359 28475
rect 35365 27673 35601 27909
rect 36237 27797 36473 28033
rect 37123 27896 37359 28132
rect 32119 27278 32355 27514
rect 32964 27350 33200 27586
rect 33720 27362 33956 27598
rect 34565 27434 34801 27670
rect 35365 27341 35601 27577
rect 36237 27465 36473 27701
rect 37123 27553 37359 27789
rect 32964 27013 33200 27249
rect 33720 27025 33956 27261
rect 34565 27097 34801 27333
rect 35365 27009 35601 27245
rect 36237 27133 36473 27369
rect 37123 27210 37359 27446
rect 37949 27413 38185 27649
rect 32964 26676 33200 26912
rect 33720 26688 33956 26924
rect 34565 26760 34801 26996
rect 35365 26677 35601 26913
rect 36237 26801 36473 27037
rect 37123 26867 37359 27103
rect 37949 27088 38185 27324
rect 37949 26763 38185 26999
rect 32964 26339 33200 26575
rect 33720 26351 33956 26587
rect 34565 26423 34801 26659
rect 35365 26344 35601 26580
rect 36237 26469 36473 26705
rect 37123 26524 37359 26760
rect 37949 26437 38185 26673
rect 38748 26614 38984 26850
rect 33720 26014 33956 26250
rect 34565 26086 34801 26322
rect 35365 26011 35601 26247
rect 36237 26137 36473 26373
rect 37123 26180 37359 26416
rect 37949 26111 38185 26347
rect 38748 26289 38984 26525
rect 33720 25677 33956 25913
rect 34565 25749 34801 25985
rect 35365 25678 35601 25914
rect 36237 25805 36473 26041
rect 37123 25836 37359 26072
rect 37949 25785 38185 26021
rect 38748 25964 38984 26200
rect 34565 25412 34801 25648
rect 35365 25345 35601 25581
rect 36237 25473 36473 25709
rect 37123 25492 37359 25728
rect 37949 25459 38185 25695
rect 38748 25639 38984 25875
rect 34565 25075 34801 25311
rect 35365 25012 35601 25248
rect 36237 25141 36473 25377
rect 37123 25148 37359 25384
rect 37949 25133 38185 25369
rect 38748 25314 38984 25550
rect 34565 24738 34801 24974
rect 35365 24679 35601 24915
rect 36237 24808 36473 25044
rect 37123 24804 37359 25040
rect 37949 24807 38185 25043
rect 38748 24989 38984 25225
rect 36237 24475 36473 24711
rect 37123 24460 37359 24696
rect 37949 24481 38185 24717
rect 38748 24663 38984 24899
rect 38748 24337 38984 24573
rect 35250 23682 35486 23918
rect 35584 23682 35820 23918
rect 35918 23682 36154 23918
rect 36252 23682 36488 23918
rect 36586 23682 36822 23918
rect 36920 23682 37156 23918
rect 37254 23682 37490 23918
rect 37588 23682 37824 23918
rect 37922 23682 38158 23918
rect 38256 23682 38492 23918
rect 38590 23682 38826 23918
rect 38924 23682 39160 23918
rect 39258 23682 39494 23918
rect 39592 23682 39828 23918
rect 35250 23360 35486 23596
rect 35584 23360 35820 23596
rect 35918 23360 36154 23596
rect 36252 23360 36488 23596
rect 36586 23360 36822 23596
rect 36920 23360 37156 23596
rect 37254 23360 37490 23596
rect 37588 23360 37824 23596
rect 37922 23360 38158 23596
rect 38256 23360 38492 23596
rect 38590 23360 38826 23596
rect 38924 23360 39160 23596
rect 39258 23360 39494 23596
rect 39592 23360 39828 23596
rect 35250 23038 35486 23274
rect 35584 23038 35820 23274
rect 35918 23038 36154 23274
rect 36252 23038 36488 23274
rect 36586 23038 36822 23274
rect 36920 23038 37156 23274
rect 37254 23038 37490 23274
rect 37588 23038 37824 23274
rect 37922 23038 38158 23274
rect 38256 23038 38492 23274
rect 38590 23038 38826 23274
rect 38924 23038 39160 23274
rect 39258 23038 39494 23274
rect 39592 23038 39828 23274
rect 35250 22716 35486 22952
rect 35584 22716 35820 22952
rect 35918 22716 36154 22952
rect 36252 22716 36488 22952
rect 36586 22716 36822 22952
rect 36920 22716 37156 22952
rect 37254 22716 37490 22952
rect 37588 22716 37824 22952
rect 37922 22716 38158 22952
rect 38256 22716 38492 22952
rect 38590 22716 38826 22952
rect 38924 22716 39160 22952
rect 39258 22716 39494 22952
rect 39592 22716 39828 22952
rect 35250 22394 35486 22630
rect 35584 22394 35820 22630
rect 35918 22394 36154 22630
rect 36252 22394 36488 22630
rect 36586 22394 36822 22630
rect 36920 22394 37156 22630
rect 37254 22394 37490 22630
rect 37588 22394 37824 22630
rect 37922 22394 38158 22630
rect 38256 22394 38492 22630
rect 38590 22394 38826 22630
rect 38924 22394 39160 22630
rect 39258 22394 39494 22630
rect 39592 22394 39828 22630
rect 35250 22072 35486 22308
rect 35584 22072 35820 22308
rect 35918 22072 36154 22308
rect 36252 22072 36488 22308
rect 36586 22072 36822 22308
rect 36920 22072 37156 22308
rect 37254 22072 37490 22308
rect 37588 22072 37824 22308
rect 37922 22072 38158 22308
rect 38256 22072 38492 22308
rect 38590 22072 38826 22308
rect 38924 22072 39160 22308
rect 39258 22072 39494 22308
rect 39592 22072 39828 22308
rect 35250 21750 35486 21986
rect 35584 21750 35820 21986
rect 35918 21750 36154 21986
rect 36252 21750 36488 21986
rect 36586 21750 36822 21986
rect 36920 21750 37156 21986
rect 37254 21750 37490 21986
rect 37588 21750 37824 21986
rect 37922 21750 38158 21986
rect 38256 21750 38492 21986
rect 38590 21750 38826 21986
rect 38924 21750 39160 21986
rect 39258 21750 39494 21986
rect 39592 21750 39828 21986
rect 35250 21428 35486 21664
rect 35584 21428 35820 21664
rect 35918 21428 36154 21664
rect 36252 21428 36488 21664
rect 36586 21428 36822 21664
rect 36920 21428 37156 21664
rect 37254 21428 37490 21664
rect 37588 21428 37824 21664
rect 37922 21428 38158 21664
rect 38256 21428 38492 21664
rect 38590 21428 38826 21664
rect 38924 21428 39160 21664
rect 39258 21428 39494 21664
rect 39592 21428 39828 21664
rect 35250 21106 35486 21342
rect 35584 21106 35820 21342
rect 35918 21106 36154 21342
rect 36252 21106 36488 21342
rect 36586 21106 36822 21342
rect 36920 21106 37156 21342
rect 37254 21106 37490 21342
rect 37588 21106 37824 21342
rect 37922 21106 38158 21342
rect 38256 21106 38492 21342
rect 38590 21106 38826 21342
rect 38924 21106 39160 21342
rect 39258 21106 39494 21342
rect 39592 21106 39828 21342
rect 35250 20784 35486 21020
rect 35584 20784 35820 21020
rect 35918 20784 36154 21020
rect 36252 20784 36488 21020
rect 36586 20784 36822 21020
rect 36920 20784 37156 21020
rect 37254 20784 37490 21020
rect 37588 20784 37824 21020
rect 37922 20784 38158 21020
rect 38256 20784 38492 21020
rect 38590 20784 38826 21020
rect 38924 20784 39160 21020
rect 39258 20784 39494 21020
rect 39592 20784 39828 21020
rect 35250 20462 35486 20698
rect 35584 20462 35820 20698
rect 35918 20462 36154 20698
rect 36252 20462 36488 20698
rect 36586 20462 36822 20698
rect 36920 20462 37156 20698
rect 37254 20462 37490 20698
rect 37588 20462 37824 20698
rect 37922 20462 38158 20698
rect 38256 20462 38492 20698
rect 38590 20462 38826 20698
rect 38924 20462 39160 20698
rect 39258 20462 39494 20698
rect 39592 20462 39828 20698
rect 35250 20140 35486 20376
rect 35584 20140 35820 20376
rect 35918 20140 36154 20376
rect 36252 20140 36488 20376
rect 36586 20140 36822 20376
rect 36920 20140 37156 20376
rect 37254 20140 37490 20376
rect 37588 20140 37824 20376
rect 37922 20140 38158 20376
rect 38256 20140 38492 20376
rect 38590 20140 38826 20376
rect 38924 20140 39160 20376
rect 39258 20140 39494 20376
rect 39592 20140 39828 20376
rect 35250 19818 35486 20054
rect 35584 19818 35820 20054
rect 35918 19818 36154 20054
rect 36252 19818 36488 20054
rect 36586 19818 36822 20054
rect 36920 19818 37156 20054
rect 37254 19818 37490 20054
rect 37588 19818 37824 20054
rect 37922 19818 38158 20054
rect 38256 19818 38492 20054
rect 38590 19818 38826 20054
rect 38924 19818 39160 20054
rect 39258 19818 39494 20054
rect 39592 19818 39828 20054
rect 529 19300 765 19536
rect 863 19300 1099 19536
rect 1197 19300 1433 19536
rect 1531 19300 1767 19536
rect 1865 19300 2101 19536
rect 2199 19300 2435 19536
rect 2533 19300 2769 19536
rect 2867 19300 3103 19536
rect 3201 19300 3437 19536
rect 3535 19300 3771 19536
rect 3869 19300 4105 19536
rect 4203 19300 4439 19536
rect 4537 19300 4773 19536
rect 4871 19300 5107 19536
rect 5205 19300 5441 19536
rect 5538 19300 5774 19536
rect 5871 19300 6107 19536
rect 6204 19300 6440 19536
rect 6537 19300 6773 19536
rect 6870 19300 7106 19536
rect 7203 19300 7439 19536
rect 7536 19300 7772 19536
rect 529 18968 765 19204
rect 863 18968 1099 19204
rect 1197 18968 1433 19204
rect 1531 18968 1767 19204
rect 1865 18968 2101 19204
rect 2199 18968 2435 19204
rect 2533 18968 2769 19204
rect 2867 18968 3103 19204
rect 3201 18968 3437 19204
rect 3535 18968 3771 19204
rect 3869 18968 4105 19204
rect 4203 18968 4439 19204
rect 4537 18968 4773 19204
rect 4871 18968 5107 19204
rect 5205 18968 5441 19204
rect 5538 18968 5774 19204
rect 5871 18968 6107 19204
rect 6204 18968 6440 19204
rect 6537 18968 6773 19204
rect 6870 18968 7106 19204
rect 7203 18968 7439 19204
rect 7536 18968 7772 19204
rect 35250 19496 35486 19732
rect 35584 19496 35820 19732
rect 35918 19496 36154 19732
rect 36252 19496 36488 19732
rect 36586 19496 36822 19732
rect 36920 19496 37156 19732
rect 37254 19496 37490 19732
rect 37588 19496 37824 19732
rect 37922 19496 38158 19732
rect 38256 19496 38492 19732
rect 38590 19496 38826 19732
rect 38924 19496 39160 19732
rect 39258 19496 39494 19732
rect 39592 19496 39828 19732
rect 35250 19174 35486 19410
rect 35584 19174 35820 19410
rect 35918 19174 36154 19410
rect 36252 19174 36488 19410
rect 36586 19174 36822 19410
rect 36920 19174 37156 19410
rect 37254 19174 37490 19410
rect 37588 19174 37824 19410
rect 37922 19174 38158 19410
rect 38256 19174 38492 19410
rect 38590 19174 38826 19410
rect 38924 19174 39160 19410
rect 39258 19174 39494 19410
rect 39592 19174 39828 19410
rect 529 18636 765 18872
rect 863 18636 1099 18872
rect 1197 18636 1433 18872
rect 1531 18636 1767 18872
rect 1865 18636 2101 18872
rect 2199 18636 2435 18872
rect 2533 18636 2769 18872
rect 2867 18636 3103 18872
rect 3201 18636 3437 18872
rect 3535 18636 3771 18872
rect 3869 18636 4105 18872
rect 4203 18636 4439 18872
rect 4537 18636 4773 18872
rect 4871 18636 5107 18872
rect 5205 18636 5441 18872
rect 5538 18636 5774 18872
rect 5871 18636 6107 18872
rect 6204 18636 6440 18872
rect 6537 18636 6773 18872
rect 6870 18636 7106 18872
rect 7203 18636 7439 18872
rect 7536 18636 7772 18872
rect 8138 18684 8374 18920
rect 529 18304 765 18540
rect 863 18304 1099 18540
rect 1197 18304 1433 18540
rect 1531 18304 1767 18540
rect 1865 18304 2101 18540
rect 2199 18304 2435 18540
rect 2533 18304 2769 18540
rect 2867 18304 3103 18540
rect 3201 18304 3437 18540
rect 3535 18304 3771 18540
rect 3869 18304 4105 18540
rect 4203 18304 4439 18540
rect 4537 18304 4773 18540
rect 4871 18304 5107 18540
rect 5205 18304 5441 18540
rect 5538 18304 5774 18540
rect 5871 18304 6107 18540
rect 6204 18304 6440 18540
rect 6537 18304 6773 18540
rect 6870 18304 7106 18540
rect 7203 18304 7439 18540
rect 7536 18304 7772 18540
rect 8138 18360 8374 18596
rect 529 17972 765 18208
rect 863 17972 1099 18208
rect 1197 17972 1433 18208
rect 1531 17972 1767 18208
rect 1865 17972 2101 18208
rect 2199 17972 2435 18208
rect 2533 17972 2769 18208
rect 2867 17972 3103 18208
rect 3201 17972 3437 18208
rect 3535 17972 3771 18208
rect 3869 17972 4105 18208
rect 4203 17972 4439 18208
rect 4537 17972 4773 18208
rect 4871 17972 5107 18208
rect 5205 17972 5441 18208
rect 5538 17972 5774 18208
rect 5871 17972 6107 18208
rect 6204 17972 6440 18208
rect 6537 17972 6773 18208
rect 6870 17972 7106 18208
rect 7203 17972 7439 18208
rect 7536 17972 7772 18208
rect 8138 18036 8374 18272
rect 35250 18852 35486 19088
rect 35584 18852 35820 19088
rect 35918 18852 36154 19088
rect 36252 18852 36488 19088
rect 36586 18852 36822 19088
rect 36920 18852 37156 19088
rect 37254 18852 37490 19088
rect 37588 18852 37824 19088
rect 37922 18852 38158 19088
rect 38256 18852 38492 19088
rect 38590 18852 38826 19088
rect 38924 18852 39160 19088
rect 39258 18852 39494 19088
rect 39592 18852 39828 19088
rect 35250 18530 35486 18766
rect 35584 18530 35820 18766
rect 35918 18530 36154 18766
rect 36252 18530 36488 18766
rect 36586 18530 36822 18766
rect 36920 18530 37156 18766
rect 37254 18530 37490 18766
rect 37588 18530 37824 18766
rect 37922 18530 38158 18766
rect 38256 18530 38492 18766
rect 38590 18530 38826 18766
rect 38924 18530 39160 18766
rect 39258 18530 39494 18766
rect 39592 18530 39828 18766
rect 8835 17987 9071 18223
rect 529 17640 765 17876
rect 863 17640 1099 17876
rect 1197 17640 1433 17876
rect 1531 17640 1767 17876
rect 1865 17640 2101 17876
rect 2199 17640 2435 17876
rect 2533 17640 2769 17876
rect 2867 17640 3103 17876
rect 3201 17640 3437 17876
rect 3535 17640 3771 17876
rect 3869 17640 4105 17876
rect 4203 17640 4439 17876
rect 4537 17640 4773 17876
rect 4871 17640 5107 17876
rect 5205 17640 5441 17876
rect 5538 17640 5774 17876
rect 5871 17640 6107 17876
rect 6204 17640 6440 17876
rect 6537 17640 6773 17876
rect 6870 17640 7106 17876
rect 7203 17640 7439 17876
rect 7536 17640 7772 17876
rect 8138 17712 8374 17948
rect 8835 17663 9071 17899
rect 529 17308 765 17544
rect 863 17308 1099 17544
rect 1197 17308 1433 17544
rect 1531 17308 1767 17544
rect 1865 17308 2101 17544
rect 2199 17308 2435 17544
rect 2533 17308 2769 17544
rect 2867 17308 3103 17544
rect 3201 17308 3437 17544
rect 3535 17308 3771 17544
rect 3869 17308 4105 17544
rect 4203 17308 4439 17544
rect 4537 17308 4773 17544
rect 4871 17308 5107 17544
rect 5205 17308 5441 17544
rect 5538 17308 5774 17544
rect 5871 17308 6107 17544
rect 6204 17308 6440 17544
rect 6537 17308 6773 17544
rect 6870 17308 7106 17544
rect 7203 17308 7439 17544
rect 7536 17308 7772 17544
rect 8138 17388 8374 17624
rect 8835 17339 9071 17575
rect 35250 18208 35486 18444
rect 35584 18208 35820 18444
rect 35918 18208 36154 18444
rect 36252 18208 36488 18444
rect 36586 18208 36822 18444
rect 36920 18208 37156 18444
rect 37254 18208 37490 18444
rect 37588 18208 37824 18444
rect 37922 18208 38158 18444
rect 38256 18208 38492 18444
rect 38590 18208 38826 18444
rect 38924 18208 39160 18444
rect 39258 18208 39494 18444
rect 39592 18208 39828 18444
rect 35250 17886 35486 18122
rect 35584 17886 35820 18122
rect 35918 17886 36154 18122
rect 36252 17886 36488 18122
rect 36586 17886 36822 18122
rect 36920 17886 37156 18122
rect 37254 17886 37490 18122
rect 37588 17886 37824 18122
rect 37922 17886 38158 18122
rect 38256 17886 38492 18122
rect 38590 17886 38826 18122
rect 38924 17886 39160 18122
rect 39258 17886 39494 18122
rect 39592 17886 39828 18122
rect 35250 17564 35486 17800
rect 35584 17564 35820 17800
rect 35918 17564 36154 17800
rect 36252 17564 36488 17800
rect 36586 17564 36822 17800
rect 36920 17564 37156 17800
rect 37254 17564 37490 17800
rect 37588 17564 37824 17800
rect 37922 17564 38158 17800
rect 38256 17564 38492 17800
rect 38590 17564 38826 17800
rect 38924 17564 39160 17800
rect 39258 17564 39494 17800
rect 39592 17564 39828 17800
rect 9494 17328 9730 17564
rect 529 16976 765 17212
rect 863 16976 1099 17212
rect 1197 16976 1433 17212
rect 1531 16976 1767 17212
rect 1865 16976 2101 17212
rect 2199 16976 2435 17212
rect 2533 16976 2769 17212
rect 2867 16976 3103 17212
rect 3201 16976 3437 17212
rect 3535 16976 3771 17212
rect 3869 16976 4105 17212
rect 4203 16976 4439 17212
rect 4537 16976 4773 17212
rect 4871 16976 5107 17212
rect 5205 16976 5441 17212
rect 5538 16976 5774 17212
rect 5871 16976 6107 17212
rect 6204 16976 6440 17212
rect 6537 16976 6773 17212
rect 6870 16976 7106 17212
rect 7203 16976 7439 17212
rect 7536 16976 7772 17212
rect 8138 17064 8374 17300
rect 8835 17015 9071 17251
rect 9494 17004 9730 17240
rect 529 16644 765 16880
rect 863 16644 1099 16880
rect 1197 16644 1433 16880
rect 1531 16644 1767 16880
rect 1865 16644 2101 16880
rect 2199 16644 2435 16880
rect 2533 16644 2769 16880
rect 2867 16644 3103 16880
rect 3201 16644 3437 16880
rect 3535 16644 3771 16880
rect 3869 16644 4105 16880
rect 4203 16644 4439 16880
rect 4537 16644 4773 16880
rect 4871 16644 5107 16880
rect 5205 16644 5441 16880
rect 5538 16644 5774 16880
rect 5871 16644 6107 16880
rect 6204 16644 6440 16880
rect 6537 16644 6773 16880
rect 6870 16644 7106 16880
rect 7203 16644 7439 16880
rect 7536 16644 7772 16880
rect 8138 16740 8374 16976
rect 8835 16691 9071 16927
rect 9494 16680 9730 16916
rect 35250 17242 35486 17478
rect 35584 17242 35820 17478
rect 35918 17242 36154 17478
rect 36252 17242 36488 17478
rect 36586 17242 36822 17478
rect 36920 17242 37156 17478
rect 37254 17242 37490 17478
rect 37588 17242 37824 17478
rect 37922 17242 38158 17478
rect 38256 17242 38492 17478
rect 38590 17242 38826 17478
rect 38924 17242 39160 17478
rect 39258 17242 39494 17478
rect 39592 17242 39828 17478
rect 35250 16920 35486 17156
rect 35584 16920 35820 17156
rect 35918 16920 36154 17156
rect 36252 16920 36488 17156
rect 36586 16920 36822 17156
rect 36920 16920 37156 17156
rect 37254 16920 37490 17156
rect 37588 16920 37824 17156
rect 37922 16920 38158 17156
rect 38256 16920 38492 17156
rect 38590 16920 38826 17156
rect 38924 16920 39160 17156
rect 39258 16920 39494 17156
rect 39592 16920 39828 17156
rect 529 16312 765 16548
rect 863 16312 1099 16548
rect 1197 16312 1433 16548
rect 1531 16312 1767 16548
rect 1865 16312 2101 16548
rect 2199 16312 2435 16548
rect 2533 16312 2769 16548
rect 2867 16312 3103 16548
rect 3201 16312 3437 16548
rect 3535 16312 3771 16548
rect 3869 16312 4105 16548
rect 4203 16312 4439 16548
rect 4537 16312 4773 16548
rect 4871 16312 5107 16548
rect 5205 16312 5441 16548
rect 5538 16312 5774 16548
rect 5871 16312 6107 16548
rect 6204 16312 6440 16548
rect 6537 16312 6773 16548
rect 6870 16312 7106 16548
rect 7203 16312 7439 16548
rect 7536 16312 7772 16548
rect 8138 16416 8374 16652
rect 10191 16631 10427 16867
rect 8835 16367 9071 16603
rect 9494 16356 9730 16592
rect 529 15980 765 16216
rect 863 15980 1099 16216
rect 1197 15980 1433 16216
rect 1531 15980 1767 16216
rect 1865 15980 2101 16216
rect 2199 15980 2435 16216
rect 2533 15980 2769 16216
rect 2867 15980 3103 16216
rect 3201 15980 3437 16216
rect 3535 15980 3771 16216
rect 3869 15980 4105 16216
rect 4203 15980 4439 16216
rect 4537 15980 4773 16216
rect 4871 15980 5107 16216
rect 5205 15980 5441 16216
rect 5538 15980 5774 16216
rect 5871 15980 6107 16216
rect 6204 15980 6440 16216
rect 6537 15980 6773 16216
rect 6870 15980 7106 16216
rect 7203 15980 7439 16216
rect 7536 15980 7772 16216
rect 8138 16092 8374 16328
rect 10191 16307 10427 16543
rect 8835 16043 9071 16279
rect 9494 16032 9730 16268
rect 529 15648 765 15884
rect 863 15648 1099 15884
rect 1197 15648 1433 15884
rect 1531 15648 1767 15884
rect 1865 15648 2101 15884
rect 2199 15648 2435 15884
rect 2533 15648 2769 15884
rect 2867 15648 3103 15884
rect 3201 15648 3437 15884
rect 3535 15648 3771 15884
rect 3869 15648 4105 15884
rect 4203 15648 4439 15884
rect 4537 15648 4773 15884
rect 4871 15648 5107 15884
rect 5205 15648 5441 15884
rect 5538 15648 5774 15884
rect 5871 15648 6107 15884
rect 6204 15648 6440 15884
rect 6537 15648 6773 15884
rect 6870 15648 7106 15884
rect 7203 15648 7439 15884
rect 7536 15648 7772 15884
rect 8138 15768 8374 16004
rect 10191 15983 10427 16219
rect 35250 16598 35486 16834
rect 35584 16598 35820 16834
rect 35918 16598 36154 16834
rect 36252 16598 36488 16834
rect 36586 16598 36822 16834
rect 36920 16598 37156 16834
rect 37254 16598 37490 16834
rect 37588 16598 37824 16834
rect 37922 16598 38158 16834
rect 38256 16598 38492 16834
rect 38590 16598 38826 16834
rect 38924 16598 39160 16834
rect 39258 16598 39494 16834
rect 39592 16598 39828 16834
rect 35250 16276 35486 16512
rect 35584 16276 35820 16512
rect 35918 16276 36154 16512
rect 36252 16276 36488 16512
rect 36586 16276 36822 16512
rect 36920 16276 37156 16512
rect 37254 16276 37490 16512
rect 37588 16276 37824 16512
rect 37922 16276 38158 16512
rect 38256 16276 38492 16512
rect 38590 16276 38826 16512
rect 38924 16276 39160 16512
rect 39258 16276 39494 16512
rect 39592 16276 39828 16512
rect 8835 15719 9071 15955
rect 10870 15952 11106 16188
rect 9494 15708 9730 15944
rect 529 15316 765 15552
rect 863 15316 1099 15552
rect 1197 15316 1433 15552
rect 1531 15316 1767 15552
rect 1865 15316 2101 15552
rect 2199 15316 2435 15552
rect 2533 15316 2769 15552
rect 2867 15316 3103 15552
rect 3201 15316 3437 15552
rect 3535 15316 3771 15552
rect 3869 15316 4105 15552
rect 4203 15316 4439 15552
rect 4537 15316 4773 15552
rect 4871 15316 5107 15552
rect 5205 15316 5441 15552
rect 5538 15316 5774 15552
rect 5871 15316 6107 15552
rect 6204 15316 6440 15552
rect 6537 15316 6773 15552
rect 6870 15316 7106 15552
rect 7203 15316 7439 15552
rect 7536 15316 7772 15552
rect 8138 15444 8374 15680
rect 10191 15659 10427 15895
rect 8835 15395 9071 15631
rect 10870 15628 11106 15864
rect 9494 15384 9730 15620
rect 529 14984 765 15220
rect 863 14984 1099 15220
rect 1197 14984 1433 15220
rect 1531 14984 1767 15220
rect 1865 14984 2101 15220
rect 2199 14984 2435 15220
rect 2533 14984 2769 15220
rect 2867 14984 3103 15220
rect 3201 14984 3437 15220
rect 3535 14984 3771 15220
rect 3869 14984 4105 15220
rect 4203 14984 4439 15220
rect 4537 14984 4773 15220
rect 4871 14984 5107 15220
rect 5205 14984 5441 15220
rect 5538 14984 5774 15220
rect 5871 14984 6107 15220
rect 6204 14984 6440 15220
rect 6537 14984 6773 15220
rect 6870 14984 7106 15220
rect 7203 14984 7439 15220
rect 7536 14984 7772 15220
rect 8138 15120 8374 15356
rect 10191 15335 10427 15571
rect 35250 15954 35486 16190
rect 35584 15954 35820 16190
rect 35918 15954 36154 16190
rect 36252 15954 36488 16190
rect 36586 15954 36822 16190
rect 36920 15954 37156 16190
rect 37254 15954 37490 16190
rect 37588 15954 37824 16190
rect 37922 15954 38158 16190
rect 38256 15954 38492 16190
rect 38590 15954 38826 16190
rect 38924 15954 39160 16190
rect 39258 15954 39494 16190
rect 39592 15954 39828 16190
rect 35250 15632 35486 15868
rect 35584 15632 35820 15868
rect 35918 15632 36154 15868
rect 36252 15632 36488 15868
rect 36586 15632 36822 15868
rect 36920 15632 37156 15868
rect 37254 15632 37490 15868
rect 37588 15632 37824 15868
rect 37922 15632 38158 15868
rect 38256 15632 38492 15868
rect 38590 15632 38826 15868
rect 38924 15632 39160 15868
rect 39258 15632 39494 15868
rect 39592 15632 39828 15868
rect 8835 15071 9071 15307
rect 10870 15304 11106 15540
rect 9494 15060 9730 15296
rect 11567 15255 11803 15491
rect 8138 14796 8374 15032
rect 10191 15011 10427 15247
rect 8835 14747 9071 14983
rect 10870 14980 11106 15216
rect 9494 14736 9730 14972
rect 11567 14931 11803 15167
rect 8138 14472 8374 14708
rect 10191 14687 10427 14923
rect 296 14154 532 14390
rect 627 14154 863 14390
rect 958 14154 1194 14390
rect 1289 14154 1525 14390
rect 1620 14154 1856 14390
rect 1951 14154 2187 14390
rect 2282 14154 2518 14390
rect 2613 14154 2849 14390
rect 2944 14154 3180 14390
rect 3275 14154 3511 14390
rect 3606 14154 3842 14390
rect 3936 14154 4172 14390
rect 4266 14154 4502 14390
rect 4596 14154 4832 14390
rect 4926 14154 5162 14390
rect 5256 14154 5492 14390
rect 8835 14423 9071 14659
rect 10870 14656 11106 14892
rect 9494 14412 9730 14648
rect 11567 14607 11803 14843
rect 35250 15310 35486 15546
rect 35584 15310 35820 15546
rect 35918 15310 36154 15546
rect 36252 15310 36488 15546
rect 36586 15310 36822 15546
rect 36920 15310 37156 15546
rect 37254 15310 37490 15546
rect 37588 15310 37824 15546
rect 37922 15310 38158 15546
rect 38256 15310 38492 15546
rect 38590 15310 38826 15546
rect 38924 15310 39160 15546
rect 39258 15310 39494 15546
rect 39592 15310 39828 15546
rect 35250 14988 35486 15224
rect 35584 14988 35820 15224
rect 35918 14988 36154 15224
rect 36252 14988 36488 15224
rect 36586 14988 36822 15224
rect 36920 14988 37156 15224
rect 37254 14988 37490 15224
rect 37588 14988 37824 15224
rect 37922 14988 38158 15224
rect 38256 14988 38492 15224
rect 38590 14988 38826 15224
rect 38924 14988 39160 15224
rect 39258 14988 39494 15224
rect 39592 14988 39828 15224
rect 8138 14148 8374 14384
rect 10191 14363 10427 14599
rect 12226 14596 12462 14832
rect 8835 14099 9071 14335
rect 10870 14332 11106 14568
rect 5581 13856 5817 14092
rect 9494 14088 9730 14324
rect 11567 14283 11803 14519
rect 296 13600 532 13836
rect 627 13600 863 13836
rect 958 13600 1194 13836
rect 1289 13600 1525 13836
rect 1620 13600 1856 13836
rect 1951 13600 2187 13836
rect 2282 13600 2518 13836
rect 2613 13600 2849 13836
rect 2944 13600 3180 13836
rect 3275 13600 3511 13836
rect 3606 13600 3842 13836
rect 3936 13600 4172 13836
rect 4266 13600 4502 13836
rect 4596 13600 4832 13836
rect 4926 13600 5162 13836
rect 5256 13600 5492 13836
rect 8138 13824 8374 14060
rect 10191 14039 10427 14275
rect 12226 14272 12462 14508
rect 8835 13775 9071 14011
rect 10870 14008 11106 14244
rect 9494 13764 9730 14000
rect 11567 13959 11803 14195
rect 5581 13309 5817 13545
rect 5985 13452 6221 13688
rect 8138 13500 8374 13736
rect 10191 13715 10427 13951
rect 12226 13948 12462 14184
rect 35250 14666 35486 14902
rect 35584 14666 35820 14902
rect 35918 14666 36154 14902
rect 36252 14666 36488 14902
rect 36586 14666 36822 14902
rect 36920 14666 37156 14902
rect 37254 14666 37490 14902
rect 37588 14666 37824 14902
rect 37922 14666 38158 14902
rect 38256 14666 38492 14902
rect 38590 14666 38826 14902
rect 38924 14666 39160 14902
rect 39258 14666 39494 14902
rect 39592 14666 39828 14902
rect 35250 14344 35486 14580
rect 35584 14344 35820 14580
rect 35918 14344 36154 14580
rect 36252 14344 36488 14580
rect 36586 14344 36822 14580
rect 36920 14344 37156 14580
rect 37254 14344 37490 14580
rect 37588 14344 37824 14580
rect 37922 14344 38158 14580
rect 38256 14344 38492 14580
rect 38590 14344 38826 14580
rect 38924 14344 39160 14580
rect 39258 14344 39494 14580
rect 39592 14344 39828 14580
rect 8835 13451 9071 13687
rect 10870 13684 11106 13920
rect 12923 13899 13159 14135
rect 9494 13440 9730 13676
rect 11567 13635 11803 13871
rect 325 12979 561 13215
rect 830 12979 1066 13215
rect 1335 12979 1571 13215
rect 1840 12979 2076 13215
rect 2345 12979 2581 13215
rect 2850 12979 3086 13215
rect 3354 12979 3590 13215
rect 3858 12979 4094 13215
rect 4362 12979 4598 13215
rect 4866 12979 5102 13215
rect 5985 12905 6221 13141
rect 6391 13046 6627 13282
rect 8138 13176 8374 13412
rect 10191 13391 10427 13627
rect 12226 13624 12462 13860
rect 8835 13127 9071 13363
rect 10870 13360 11106 13596
rect 12923 13575 13159 13811
rect 9494 13116 9730 13352
rect 11567 13311 11803 13547
rect 325 12441 561 12677
rect 830 12441 1066 12677
rect 1335 12441 1571 12677
rect 1840 12441 2076 12677
rect 2345 12441 2581 12677
rect 2850 12441 3086 12677
rect 3354 12441 3590 12677
rect 3858 12441 4094 12677
rect 4362 12441 4598 12677
rect 4866 12441 5102 12677
rect 5220 12606 5456 12842
rect 5220 12059 5456 12295
rect 5581 12242 5817 12478
rect 6391 12499 6627 12735
rect 6795 12642 7031 12878
rect 8138 12852 8374 13088
rect 10191 13067 10427 13303
rect 12226 13300 12462 13536
rect 35250 14022 35486 14258
rect 35584 14022 35820 14258
rect 35918 14022 36154 14258
rect 36252 14022 36488 14258
rect 36586 14022 36822 14258
rect 36920 14022 37156 14258
rect 37254 14022 37490 14258
rect 37588 14022 37824 14258
rect 37922 14022 38158 14258
rect 38256 14022 38492 14258
rect 38590 14022 38826 14258
rect 38924 14022 39160 14258
rect 39258 14022 39494 14258
rect 39592 14022 39828 14258
rect 35250 13700 35486 13936
rect 35584 13700 35820 13936
rect 35918 13700 36154 13936
rect 36252 13700 36488 13936
rect 36586 13700 36822 13936
rect 36920 13700 37156 13936
rect 37254 13700 37490 13936
rect 37588 13700 37824 13936
rect 37922 13700 38158 13936
rect 38256 13700 38492 13936
rect 38590 13700 38826 13936
rect 38924 13700 39160 13936
rect 39258 13700 39494 13936
rect 39592 13700 39828 13936
rect 8835 12803 9071 13039
rect 10870 13036 11106 13272
rect 12923 13251 13159 13487
rect 13547 13275 13783 13511
rect 9494 12792 9730 13028
rect 11567 12987 11803 13223
rect 8138 12527 8374 12763
rect 10191 12743 10427 12979
rect 12226 12976 12462 13212
rect 8835 12479 9071 12715
rect 10870 12712 11106 12948
rect 12923 12927 13159 13163
rect 13547 12951 13783 13187
rect 5581 11695 5817 11931
rect 5985 11838 6221 12074
rect 6795 12095 7031 12331
rect 7194 12243 7430 12479
rect 9494 12468 9730 12704
rect 11567 12663 11803 12899
rect 10191 12419 10427 12655
rect 12226 12652 12462 12888
rect 8835 12155 9071 12391
rect 10870 12388 11106 12624
rect 12923 12603 13159 12839
rect 13547 12627 13783 12863
rect 35250 13378 35486 13614
rect 35584 13378 35820 13614
rect 35918 13378 36154 13614
rect 36252 13378 36488 13614
rect 36586 13378 36822 13614
rect 36920 13378 37156 13614
rect 37254 13378 37490 13614
rect 37588 13378 37824 13614
rect 37922 13378 38158 13614
rect 38256 13378 38492 13614
rect 38590 13378 38826 13614
rect 38924 13378 39160 13614
rect 39258 13378 39494 13614
rect 39592 13378 39828 13614
rect 35250 13056 35486 13292
rect 35584 13056 35820 13292
rect 35918 13056 36154 13292
rect 36252 13056 36488 13292
rect 36586 13056 36822 13292
rect 36920 13056 37156 13292
rect 37254 13056 37490 13292
rect 37588 13056 37824 13292
rect 37922 13056 38158 13292
rect 38256 13056 38492 13292
rect 38590 13056 38826 13292
rect 38924 13056 39160 13292
rect 39258 13056 39494 13292
rect 39592 13056 39828 13292
rect 14244 12578 14480 12814
rect 9494 12144 9730 12380
rect 11567 12339 11803 12575
rect 10191 12095 10427 12331
rect 12226 12328 12462 12564
rect 7194 11696 7430 11932
rect 7598 11839 7834 12075
rect 8835 11830 9071 12066
rect 10870 12064 11106 12300
rect 12923 12279 13159 12515
rect 13547 12303 13783 12539
rect 14244 12256 14480 12492
rect 9494 11820 9730 12056
rect 11567 12015 11803 12251
rect 5985 11291 6221 11527
rect 6391 11432 6627 11668
rect 6391 10885 6627 11121
rect 6800 11026 7036 11262
rect 7598 11292 7834 11528
rect 8009 11428 8245 11664
rect 10191 11771 10427 12007
rect 12226 12004 12462 12240
rect 10870 11740 11106 11976
rect 12923 11955 13159 12191
rect 13547 11979 13783 12215
rect 14244 11934 14480 12170
rect 35250 12734 35486 12970
rect 35584 12734 35820 12970
rect 35918 12734 36154 12970
rect 36252 12734 36488 12970
rect 36586 12734 36822 12970
rect 36920 12734 37156 12970
rect 37254 12734 37490 12970
rect 37588 12734 37824 12970
rect 37922 12734 38158 12970
rect 38256 12734 38492 12970
rect 38590 12734 38826 12970
rect 38924 12734 39160 12970
rect 39258 12734 39494 12970
rect 39592 12734 39828 12970
rect 35250 12412 35486 12648
rect 35584 12412 35820 12648
rect 35918 12412 36154 12648
rect 36252 12412 36488 12648
rect 36586 12412 36822 12648
rect 36920 12412 37156 12648
rect 37254 12412 37490 12648
rect 37588 12412 37824 12648
rect 37922 12412 38158 12648
rect 38256 12412 38492 12648
rect 38590 12412 38826 12648
rect 38924 12412 39160 12648
rect 39258 12412 39494 12648
rect 39592 12412 39828 12648
rect 9494 11496 9730 11732
rect 11567 11691 11803 11927
rect 14903 11919 15139 12155
rect 10191 11447 10427 11683
rect 12226 11680 12462 11916
rect 10870 11416 11106 11652
rect 12923 11631 13159 11867
rect 13547 11655 13783 11891
rect 14244 11612 14480 11848
rect 6800 10479 7036 10715
rect 7161 10662 7397 10898
rect 8009 10881 8245 11117
rect 8413 11024 8649 11260
rect 9494 11171 9730 11407
rect 11567 11367 11803 11603
rect 14903 11598 15139 11834
rect 10191 11123 10427 11359
rect 12226 11356 12462 11592
rect 10870 11092 11106 11328
rect 12923 11307 13159 11543
rect 13547 11331 13783 11567
rect 14244 11290 14480 11526
rect 11567 11043 11803 11279
rect 14903 11277 15139 11513
rect 35250 12090 35486 12326
rect 35584 12090 35820 12326
rect 35918 12090 36154 12326
rect 36252 12090 36488 12326
rect 36586 12090 36822 12326
rect 36920 12090 37156 12326
rect 37254 12090 37490 12326
rect 37588 12090 37824 12326
rect 37922 12090 38158 12326
rect 38256 12090 38492 12326
rect 38590 12090 38826 12326
rect 38924 12090 39160 12326
rect 39258 12090 39494 12326
rect 39592 12090 39828 12326
rect 35250 11768 35486 12004
rect 35584 11768 35820 12004
rect 35918 11768 36154 12004
rect 36252 11768 36488 12004
rect 36586 11768 36822 12004
rect 36920 11768 37156 12004
rect 37254 11768 37490 12004
rect 37588 11768 37824 12004
rect 37922 11768 38158 12004
rect 38256 11768 38492 12004
rect 38590 11768 38826 12004
rect 38924 11768 39160 12004
rect 39258 11768 39494 12004
rect 39592 11768 39828 12004
rect 7161 10115 7397 10351
rect 7565 10258 7801 10494
rect 8413 10477 8649 10713
rect 8812 10625 9048 10861
rect 10191 10799 10427 11035
rect 12226 11032 12462 11268
rect 10870 10768 11106 11004
rect 12923 10983 13159 11219
rect 13547 11007 13783 11243
rect 15600 11222 15836 11458
rect 14244 10968 14480 11204
rect 14903 10956 15139 11192
rect 11567 10719 11803 10955
rect 295 9684 531 9920
rect 830 9684 1066 9920
rect 1365 9684 1601 9920
rect 1900 9684 2136 9920
rect 2434 9684 2670 9920
rect 2968 9684 3204 9920
rect 3502 9684 3738 9920
rect 7565 9711 7801 9947
rect 7971 9852 8207 10088
rect 8812 10078 9048 10314
rect 9216 10221 9452 10457
rect 10191 10474 10427 10710
rect 12226 10708 12462 10944
rect 10870 10444 11106 10680
rect 12923 10659 13159 10895
rect 13547 10683 13783 10919
rect 15600 10891 15836 11127
rect 35250 11446 35486 11682
rect 35584 11446 35820 11682
rect 35918 11446 36154 11682
rect 36252 11446 36488 11682
rect 36586 11446 36822 11682
rect 36920 11446 37156 11682
rect 37254 11446 37490 11682
rect 37588 11446 37824 11682
rect 37922 11446 38158 11682
rect 38256 11446 38492 11682
rect 38590 11446 38826 11682
rect 38924 11446 39160 11682
rect 39258 11446 39494 11682
rect 39592 11446 39828 11682
rect 35250 11124 35486 11360
rect 35584 11124 35820 11360
rect 35918 11124 36154 11360
rect 36252 11124 36488 11360
rect 36586 11124 36822 11360
rect 36920 11124 37156 11360
rect 37254 11124 37490 11360
rect 37588 11124 37824 11360
rect 37922 11124 38158 11360
rect 38256 11124 38492 11360
rect 38590 11124 38826 11360
rect 38924 11124 39160 11360
rect 39258 11124 39494 11360
rect 39592 11124 39828 11360
rect 14244 10646 14480 10882
rect 14903 10635 15139 10871
rect 16073 10861 16309 11097
rect 11567 10395 11803 10631
rect 12226 10384 12462 10620
rect 295 9110 531 9346
rect 830 9110 1066 9346
rect 1365 9110 1601 9346
rect 1900 9110 2136 9346
rect 2434 9110 2670 9346
rect 2968 9110 3204 9346
rect 3502 9110 3738 9346
rect 3820 9305 4056 9541
rect 7971 9305 8207 9541
rect 8365 9461 8601 9697
rect 9216 9674 9452 9910
rect 9649 9788 9885 10024
rect 10870 10120 11106 10356
rect 12923 10335 13159 10571
rect 13547 10359 13783 10595
rect 15600 10560 15836 10796
rect 14244 10324 14480 10560
rect 14903 10314 15139 10550
rect 11567 10071 11803 10307
rect 12226 10060 12462 10296
rect 10870 9795 11106 10031
rect 12923 10011 13159 10247
rect 13547 10035 13783 10271
rect 14244 10002 14480 10238
rect 15600 10229 15836 10465
rect 14903 9993 15139 10229
rect 16073 10226 16309 10462
rect 35250 10802 35486 11038
rect 35584 10802 35820 11038
rect 35918 10802 36154 11038
rect 36252 10802 36488 11038
rect 36586 10802 36822 11038
rect 36920 10802 37156 11038
rect 37254 10802 37490 11038
rect 37588 10802 37824 11038
rect 37922 10802 38158 11038
rect 38256 10802 38492 11038
rect 38590 10802 38826 11038
rect 38924 10802 39160 11038
rect 39258 10802 39494 11038
rect 39592 10802 39828 11038
rect 35250 10480 35486 10716
rect 35584 10480 35820 10716
rect 35918 10480 36154 10716
rect 36252 10480 36488 10716
rect 36586 10480 36822 10716
rect 36920 10480 37156 10716
rect 37254 10480 37490 10716
rect 37588 10480 37824 10716
rect 37922 10480 38158 10716
rect 38256 10480 38492 10716
rect 38590 10480 38826 10716
rect 38924 10480 39160 10716
rect 39258 10480 39494 10716
rect 39592 10480 39828 10716
rect 11567 9747 11803 9983
rect 12226 9736 12462 9972
rect 12923 9687 13159 9923
rect 13547 9711 13783 9947
rect 14244 9679 14480 9915
rect 14903 9672 15139 9908
rect 15600 9898 15836 10134
rect 16050 9843 16286 10079
rect 16545 9843 16781 10079
rect 17039 9843 17275 10079
rect 267 8466 503 8702
rect 816 8466 1052 8702
rect 1365 8466 1601 8702
rect 1914 8466 2150 8702
rect 2463 8466 2699 8702
rect 3012 8466 3248 8702
rect 3820 8758 4056 8994
rect 4195 8946 4431 9182
rect 8365 8914 8601 9150
rect 8726 9097 8962 9333
rect 9649 9241 9885 9477
rect 10053 9384 10289 9620
rect 11567 9423 11803 9659
rect 12226 9412 12462 9648
rect 12923 9363 13159 9599
rect 13547 9387 13783 9623
rect 14244 9356 14480 9592
rect 14903 9351 15139 9587
rect 15600 9567 15836 9803
rect 35250 10158 35486 10394
rect 35584 10158 35820 10394
rect 35918 10158 36154 10394
rect 36252 10158 36488 10394
rect 36586 10158 36822 10394
rect 36920 10158 37156 10394
rect 37254 10158 37490 10394
rect 37588 10158 37824 10394
rect 37922 10158 38158 10394
rect 38256 10158 38492 10394
rect 38590 10158 38826 10394
rect 38924 10158 39160 10394
rect 39258 10158 39494 10394
rect 39592 10158 39828 10394
rect 35250 9836 35486 10072
rect 35584 9836 35820 10072
rect 35918 9836 36154 10072
rect 36252 9836 36488 10072
rect 36586 9836 36822 10072
rect 36920 9836 37156 10072
rect 37254 9836 37490 10072
rect 37588 9836 37824 10072
rect 37922 9836 38158 10072
rect 38256 9836 38492 10072
rect 38590 9836 38826 10072
rect 38924 9836 39160 10072
rect 39258 9836 39494 10072
rect 39592 9836 39828 10072
rect 267 8126 503 8362
rect 816 8126 1052 8362
rect 1365 8126 1601 8362
rect 1914 8126 2150 8362
rect 2463 8126 2699 8362
rect 3012 8126 3248 8362
rect 4195 8399 4431 8635
rect 4556 8582 4792 8818
rect 8726 8550 8962 8786
rect 9130 8693 9366 8929
rect 10053 8837 10289 9073
rect 10452 8985 10688 9221
rect 11567 9098 11803 9334
rect 12226 9088 12462 9324
rect 12923 9039 13159 9275
rect 13547 9063 13783 9299
rect 14244 9033 14480 9269
rect 14903 9030 15139 9266
rect 15600 9235 15836 9471
rect 16065 9363 16301 9599
rect 16575 9363 16811 9599
rect 17084 9363 17320 9599
rect 17593 9363 17829 9599
rect 4556 8035 4792 8271
rect 4945 8196 5181 8432
rect 277 7502 513 7738
rect 860 7502 1096 7738
rect 1442 7502 1678 7738
rect 2024 7502 2260 7738
rect 2606 7502 2842 7738
rect 277 7164 513 7400
rect 860 7164 1096 7400
rect 1442 7164 1678 7400
rect 2024 7164 2260 7400
rect 2606 7164 2842 7400
rect 4945 7649 5181 7885
rect 5306 7832 5542 8068
rect 9130 8146 9366 8382
rect 9536 8287 9772 8523
rect 10452 8438 10688 8674
rect 10856 8581 11092 8817
rect 12226 8764 12462 9000
rect 12923 8715 13159 8951
rect 13547 8739 13783 8975
rect 14244 8710 14480 8946
rect 14903 8709 15139 8945
rect 15600 8903 15836 9139
rect 16065 9025 16301 9261
rect 16575 9025 16811 9261
rect 17084 9025 17320 9261
rect 17593 9025 17829 9261
rect 5306 7285 5542 7521
rect 5692 7433 5928 7669
rect 9536 7740 9772 7976
rect 9955 7871 10191 8107
rect 10856 8034 11092 8270
rect 11303 8134 11539 8370
rect 12226 8439 12462 8675
rect 12923 8391 13159 8627
rect 13547 8415 13783 8651
rect 14244 8387 14480 8623
rect 14903 8388 15139 8624
rect 15600 8571 15836 8807
rect 16065 8687 16301 8923
rect 16575 8687 16811 8923
rect 17084 8687 17320 8923
rect 17593 8687 17829 8923
rect 35250 9514 35486 9750
rect 35584 9514 35820 9750
rect 35918 9514 36154 9750
rect 36252 9514 36488 9750
rect 36586 9514 36822 9750
rect 36920 9514 37156 9750
rect 37254 9514 37490 9750
rect 37588 9514 37824 9750
rect 37922 9514 38158 9750
rect 38256 9514 38492 9750
rect 38590 9514 38826 9750
rect 38924 9514 39160 9750
rect 39258 9514 39494 9750
rect 39592 9514 39828 9750
rect 35250 9192 35486 9428
rect 35584 9192 35820 9428
rect 35918 9192 36154 9428
rect 36252 9192 36488 9428
rect 36586 9192 36822 9428
rect 36920 9192 37156 9428
rect 37254 9192 37490 9428
rect 37588 9192 37824 9428
rect 37922 9192 38158 9428
rect 38256 9192 38492 9428
rect 38590 9192 38826 9428
rect 38924 9192 39160 9428
rect 39258 9192 39494 9428
rect 39592 9192 39828 9428
rect 35250 8870 35486 9106
rect 35584 8870 35820 9106
rect 35918 8870 36154 9106
rect 36252 8870 36488 9106
rect 36586 8870 36822 9106
rect 36920 8870 37156 9106
rect 37254 8870 37490 9106
rect 37588 8870 37824 9106
rect 37922 8870 38158 9106
rect 38256 8870 38492 9106
rect 38590 8870 38826 9106
rect 38924 8870 39160 9106
rect 39258 8870 39494 9106
rect 39592 8870 39828 9106
rect 35250 8548 35486 8784
rect 35584 8548 35820 8784
rect 35918 8548 36154 8784
rect 36252 8548 36488 8784
rect 36586 8548 36822 8784
rect 36920 8548 37156 8784
rect 37254 8548 37490 8784
rect 37588 8548 37824 8784
rect 37922 8548 38158 8784
rect 38256 8548 38492 8784
rect 38590 8548 38826 8784
rect 38924 8548 39160 8784
rect 39258 8548 39494 8784
rect 39592 8548 39828 8784
rect 12923 8067 13159 8303
rect 13547 8091 13783 8327
rect 14244 8064 14480 8300
rect 14903 8066 15139 8302
rect 15600 8239 15836 8475
rect 16047 8265 16283 8501
rect 16549 8265 16785 8501
rect 17050 8265 17286 8501
rect 17551 8265 17787 8501
rect 18052 8265 18288 8501
rect 18553 8265 18789 8501
rect 5692 6886 5928 7122
rect 6067 7074 6303 7310
rect 9955 7324 10191 7560
rect 10316 7507 10552 7743
rect 11303 7587 11539 7823
rect 11707 7730 11943 7966
rect 12923 7742 13159 7978
rect 13547 7767 13783 8003
rect 14244 7741 14480 7977
rect 14903 7744 15139 7980
rect 15600 7907 15836 8143
rect 16047 7853 16283 8089
rect 16549 7853 16785 8089
rect 17050 7853 17286 8089
rect 17551 7853 17787 8089
rect 18052 7853 18288 8089
rect 18553 7853 18789 8089
rect 320 6513 556 6749
rect 786 6513 1022 6749
rect 1252 6513 1488 6749
rect 1718 6513 1954 6749
rect 2183 6513 2419 6749
rect 2506 6235 2742 6471
rect 320 5979 556 6215
rect 786 5979 1022 6215
rect 1252 5979 1488 6215
rect 1718 5979 1954 6215
rect 2183 5979 2419 6215
rect 2506 5908 2742 6144
rect 6067 6527 6303 6763
rect 6428 6710 6664 6946
rect 10316 6960 10552 7196
rect 10720 7103 10956 7339
rect 11707 7183 11943 7419
rect 12106 7331 12342 7567
rect 13547 7443 13783 7679
rect 14244 7418 14480 7654
rect 14903 7422 15139 7658
rect 15600 7575 15836 7811
rect 2888 5853 3124 6089
rect 6428 6163 6664 6399
rect 6817 6324 7053 6560
rect 10720 6556 10956 6792
rect 11126 6697 11362 6933
rect 12106 6784 12342 7020
rect 12510 6927 12746 7163
rect 13547 7118 13783 7354
rect 14244 7095 14480 7331
rect 14903 7100 15139 7336
rect 15600 7243 15836 7479
rect 16047 7441 16283 7677
rect 16549 7441 16785 7677
rect 17050 7441 17286 7677
rect 17551 7441 17787 7677
rect 18052 7441 18288 7677
rect 18553 7441 18789 7677
rect 15600 6911 15836 7147
rect 16047 7029 16283 7265
rect 16549 7029 16785 7265
rect 17050 7029 17286 7265
rect 17551 7029 17787 7265
rect 18052 7029 18288 7265
rect 18553 7029 18789 7265
rect 305 5306 541 5542
rect 772 5306 1008 5542
rect 1239 5306 1475 5542
rect 1706 5306 1942 5542
rect 2506 5580 2742 5816
rect 2888 5526 3124 5762
rect 3301 5440 3537 5676
rect 6817 5777 7053 6013
rect 7178 5960 7414 6196
rect 11126 6150 11362 6386
rect 12510 6380 12746 6616
rect 16047 6617 16283 6853
rect 16549 6617 16785 6853
rect 17050 6617 17286 6853
rect 17551 6617 17787 6853
rect 18052 6617 18288 6853
rect 18553 6617 18789 6853
rect 12869 6043 13105 6279
rect 13421 6043 13657 6279
rect 2888 5198 3124 5434
rect 305 4744 541 4980
rect 772 4744 1008 4980
rect 1239 4744 1475 4980
rect 1706 4744 1942 4980
rect 2139 4885 2375 5121
rect 3301 5113 3537 5349
rect 2139 4558 2375 4794
rect 3683 5058 3919 5294
rect 7178 5413 7414 5649
rect 7589 5552 7825 5788
rect 11703 5576 11939 5812
rect 12237 5576 12473 5812
rect 3301 4785 3537 5021
rect 2521 4503 2757 4739
rect 3683 4731 3919 4967
rect 7589 5005 7825 5241
rect 7950 5188 8186 5424
rect 294 4097 530 4333
rect 747 4097 983 4333
rect 1200 4097 1436 4333
rect 2139 4230 2375 4466
rect 2521 4176 2757 4412
rect 3683 4403 3919 4639
rect 4131 4610 4367 4846
rect 7950 4641 8186 4877
rect 2867 4157 3103 4393
rect 4131 4283 4367 4519
rect 4513 4228 4749 4464
rect 294 3769 530 4005
rect 747 3769 983 4005
rect 1200 3769 1436 4005
rect 2521 3848 2757 4084
rect 2867 3830 3103 4066
rect 3249 3775 3485 4011
rect 2867 3502 3103 3738
rect 3249 3448 3485 3684
rect 4131 3955 4367 4191
rect 4513 3901 4749 4137
rect 8366 4219 8602 4455
rect 8956 4219 9192 4455
rect 4911 3830 5147 4066
rect 757 3126 993 3362
rect 3628 3396 3864 3632
rect 4513 3573 4749 3809
rect 4911 3503 5147 3739
rect 3249 3120 3485 3356
rect 3628 3069 3864 3305
rect 4911 3175 5147 3411
rect 7402 3726 7638 3962
rect 7750 3726 7986 3962
rect 6428 3320 6664 3556
rect 6782 3320 7018 3556
rect 757 2513 993 2749
rect 1151 2732 1387 2968
rect 3628 2741 3864 2977
rect 5233 2910 5469 3146
rect 5787 2910 6023 3146
rect 1496 2387 1732 2623
rect 1151 2119 1387 2355
rect 4011 2395 4247 2631
rect 4597 2395 4833 2631
rect 1496 1774 1732 2010
rect 1836 1485 2072 1721
rect 2416 1485 2652 1721
rect 470 989 706 1225
rect 834 989 1070 1225
rect 1198 989 1434 1225
rect 470 513 706 749
rect 834 513 1070 749
rect 1198 513 1434 749
rect 470 36 706 272
rect 834 36 1070 272
rect 1198 36 1434 272
rect 1836 1122 2072 1358
rect 2416 1122 2652 1358
rect 1836 759 2072 995
rect 2416 759 2652 995
rect 1836 395 2072 631
rect 2416 395 2652 631
rect 1836 31 2072 267
rect 2416 31 2652 267
rect 3037 1893 3273 2129
rect 3393 1893 3629 2129
rect 3037 1522 3273 1758
rect 3393 1522 3629 1758
rect 3037 1151 3273 1387
rect 3393 1151 3629 1387
rect 3037 779 3273 1015
rect 3393 779 3629 1015
rect 3037 407 3273 643
rect 3393 407 3629 643
rect 3037 35 3273 271
rect 3393 35 3629 271
rect 4011 2059 4247 2295
rect 4597 2059 4833 2295
rect 4011 1723 4247 1959
rect 4597 1723 4833 1959
rect 4011 1387 4247 1623
rect 4597 1387 4833 1623
rect 4011 1051 4247 1287
rect 4597 1051 4833 1287
rect 4011 715 4247 951
rect 4597 715 4833 951
rect 4011 379 4247 615
rect 4597 379 4833 615
rect 4011 43 4247 279
rect 4597 43 4833 279
rect 5233 2551 5469 2787
rect 5787 2551 6023 2787
rect 5233 2192 5469 2428
rect 5787 2192 6023 2428
rect 5233 1833 5469 2069
rect 5787 1833 6023 2069
rect 5233 1474 5469 1710
rect 5787 1474 6023 1710
rect 5233 1114 5469 1350
rect 5787 1114 6023 1350
rect 5233 754 5469 990
rect 5787 754 6023 990
rect 5233 394 5469 630
rect 5787 394 6023 630
rect 5233 34 5469 270
rect 5787 34 6023 270
rect 6428 2992 6664 3228
rect 6782 2992 7018 3228
rect 6428 2664 6664 2900
rect 6782 2664 7018 2900
rect 6428 2336 6664 2572
rect 6782 2336 7018 2572
rect 6428 2008 6664 2244
rect 6782 2008 7018 2244
rect 6428 1680 6664 1916
rect 6782 1680 7018 1916
rect 6428 1352 6664 1588
rect 6782 1352 7018 1588
rect 6428 1024 6664 1260
rect 6782 1024 7018 1260
rect 6428 695 6664 931
rect 6782 695 7018 931
rect 6428 366 6664 602
rect 6782 366 7018 602
rect 6428 37 6664 273
rect 6782 37 7018 273
rect 7402 3397 7638 3633
rect 7750 3397 7986 3633
rect 7402 3068 7638 3304
rect 7750 3068 7986 3304
rect 7402 2739 7638 2975
rect 7750 2739 7986 2975
rect 7402 2410 7638 2646
rect 7750 2410 7986 2646
rect 7402 2081 7638 2317
rect 7750 2081 7986 2317
rect 7402 1752 7638 1988
rect 7750 1752 7986 1988
rect 7402 1423 7638 1659
rect 7750 1423 7986 1659
rect 7402 1093 7638 1329
rect 7750 1093 7986 1329
rect 7402 763 7638 999
rect 7750 763 7986 999
rect 7402 433 7638 669
rect 7750 433 7986 669
rect 7402 103 7638 339
rect 7750 103 7986 339
rect 8366 3898 8602 4134
rect 8956 3898 9192 4134
rect 8366 3577 8602 3813
rect 8956 3577 9192 3813
rect 8366 3256 8602 3492
rect 8956 3256 9192 3492
rect 8366 2935 8602 3171
rect 8956 2935 9192 3171
rect 8366 2613 8602 2849
rect 8956 2613 9192 2849
rect 8366 2291 8602 2527
rect 8956 2291 9192 2527
rect 8366 1969 8602 2205
rect 8956 1969 9192 2205
rect 8366 1647 8602 1883
rect 8956 1647 9192 1883
rect 8366 1325 8602 1561
rect 8956 1325 9192 1561
rect 8366 1003 8602 1239
rect 8956 1003 9192 1239
rect 8366 681 8602 917
rect 8956 681 9192 917
rect 8366 359 8602 595
rect 8956 359 9192 595
rect 8366 37 8602 273
rect 8956 37 9192 273
rect 11703 5251 11939 5487
rect 12237 5251 12473 5487
rect 11703 4926 11939 5162
rect 12237 4926 12473 5162
rect 11703 4601 11939 4837
rect 12237 4601 12473 4837
rect 11703 4276 11939 4512
rect 12237 4276 12473 4512
rect 11703 3951 11939 4187
rect 12237 3951 12473 4187
rect 11703 3626 11939 3862
rect 12237 3626 12473 3862
rect 11703 3301 11939 3537
rect 12237 3301 12473 3537
rect 11703 2975 11939 3211
rect 12237 2975 12473 3211
rect 11703 2649 11939 2885
rect 12237 2649 12473 2885
rect 11703 2323 11939 2559
rect 12237 2323 12473 2559
rect 11703 1997 11939 2233
rect 12237 1997 12473 2233
rect 11703 1671 11939 1907
rect 12237 1671 12473 1907
rect 11703 1345 11939 1581
rect 12237 1345 12473 1581
rect 11703 1019 11939 1255
rect 12237 1019 12473 1255
rect 11703 693 11939 929
rect 12237 693 12473 929
rect 11703 367 11939 603
rect 12237 367 12473 603
rect 11703 41 11939 277
rect 12237 41 12473 277
rect 12869 5712 13105 5948
rect 13421 5712 13657 5948
rect 12869 5381 13105 5617
rect 13421 5381 13657 5617
rect 12869 5050 13105 5286
rect 13421 5050 13657 5286
rect 12869 4719 13105 4955
rect 13421 4719 13657 4955
rect 12869 4388 13105 4624
rect 13421 4388 13657 4624
rect 12869 4057 13105 4293
rect 13421 4057 13657 4293
rect 12869 3726 13105 3962
rect 13421 3726 13657 3962
rect 12869 3395 13105 3631
rect 13421 3395 13657 3631
rect 12869 3064 13105 3300
rect 13421 3064 13657 3300
rect 12869 2733 13105 2969
rect 13421 2733 13657 2969
rect 12869 2402 13105 2638
rect 13421 2402 13657 2638
rect 12869 2071 13105 2307
rect 13421 2071 13657 2307
rect 12869 1740 13105 1976
rect 13421 1740 13657 1976
rect 12869 1408 13105 1644
rect 13421 1408 13657 1644
rect 12869 1076 13105 1312
rect 13421 1076 13657 1312
rect 12869 744 13105 980
rect 13421 744 13657 980
rect 12869 412 13105 648
rect 13421 412 13657 648
rect 12869 80 13105 316
rect 13421 80 13657 316
rect 14300 6253 14536 6489
rect 14624 6253 14860 6489
rect 14948 6253 15184 6489
rect 15272 6253 15508 6489
rect 15596 6253 15832 6489
rect 15920 6253 16156 6489
rect 16244 6253 16480 6489
rect 16568 6253 16804 6489
rect 16892 6253 17128 6489
rect 17216 6253 17452 6489
rect 17540 6253 17776 6489
rect 17864 6253 18100 6489
rect 18188 6253 18424 6489
rect 18512 6253 18748 6489
rect 14300 5923 14536 6159
rect 14624 5923 14860 6159
rect 14948 5923 15184 6159
rect 15272 5923 15508 6159
rect 15596 5923 15832 6159
rect 15920 5923 16156 6159
rect 16244 5923 16480 6159
rect 16568 5923 16804 6159
rect 16892 5923 17128 6159
rect 17216 5923 17452 6159
rect 17540 5923 17776 6159
rect 17864 5923 18100 6159
rect 18188 5923 18424 6159
rect 18512 5923 18748 6159
rect 14300 5593 14536 5829
rect 14624 5593 14860 5829
rect 14948 5593 15184 5829
rect 15272 5593 15508 5829
rect 15596 5593 15832 5829
rect 15920 5593 16156 5829
rect 16244 5593 16480 5829
rect 16568 5593 16804 5829
rect 16892 5593 17128 5829
rect 17216 5593 17452 5829
rect 17540 5593 17776 5829
rect 17864 5593 18100 5829
rect 18188 5593 18424 5829
rect 18512 5593 18748 5829
rect 14300 5263 14536 5499
rect 14624 5263 14860 5499
rect 14948 5263 15184 5499
rect 15272 5263 15508 5499
rect 15596 5263 15832 5499
rect 15920 5263 16156 5499
rect 16244 5263 16480 5499
rect 16568 5263 16804 5499
rect 16892 5263 17128 5499
rect 17216 5263 17452 5499
rect 17540 5263 17776 5499
rect 17864 5263 18100 5499
rect 18188 5263 18424 5499
rect 18512 5263 18748 5499
rect 14300 4933 14536 5169
rect 14624 4933 14860 5169
rect 14948 4933 15184 5169
rect 15272 4933 15508 5169
rect 15596 4933 15832 5169
rect 15920 4933 16156 5169
rect 16244 4933 16480 5169
rect 16568 4933 16804 5169
rect 16892 4933 17128 5169
rect 17216 4933 17452 5169
rect 17540 4933 17776 5169
rect 17864 4933 18100 5169
rect 18188 4933 18424 5169
rect 18512 4933 18748 5169
rect 14300 4603 14536 4839
rect 14624 4603 14860 4839
rect 14948 4603 15184 4839
rect 15272 4603 15508 4839
rect 15596 4603 15832 4839
rect 15920 4603 16156 4839
rect 16244 4603 16480 4839
rect 16568 4603 16804 4839
rect 16892 4603 17128 4839
rect 17216 4603 17452 4839
rect 17540 4603 17776 4839
rect 17864 4603 18100 4839
rect 18188 4603 18424 4839
rect 18512 4603 18748 4839
rect 14300 4273 14536 4509
rect 14624 4273 14860 4509
rect 14948 4273 15184 4509
rect 15272 4273 15508 4509
rect 15596 4273 15832 4509
rect 15920 4273 16156 4509
rect 16244 4273 16480 4509
rect 16568 4273 16804 4509
rect 16892 4273 17128 4509
rect 17216 4273 17452 4509
rect 17540 4273 17776 4509
rect 17864 4273 18100 4509
rect 18188 4273 18424 4509
rect 18512 4273 18748 4509
rect 14300 3943 14536 4179
rect 14624 3943 14860 4179
rect 14948 3943 15184 4179
rect 15272 3943 15508 4179
rect 15596 3943 15832 4179
rect 15920 3943 16156 4179
rect 16244 3943 16480 4179
rect 16568 3943 16804 4179
rect 16892 3943 17128 4179
rect 17216 3943 17452 4179
rect 17540 3943 17776 4179
rect 17864 3943 18100 4179
rect 18188 3943 18424 4179
rect 18512 3943 18748 4179
rect 14300 3613 14536 3849
rect 14624 3613 14860 3849
rect 14948 3613 15184 3849
rect 15272 3613 15508 3849
rect 15596 3613 15832 3849
rect 15920 3613 16156 3849
rect 16244 3613 16480 3849
rect 16568 3613 16804 3849
rect 16892 3613 17128 3849
rect 17216 3613 17452 3849
rect 17540 3613 17776 3849
rect 17864 3613 18100 3849
rect 18188 3613 18424 3849
rect 18512 3613 18748 3849
rect 14300 3283 14536 3519
rect 14624 3283 14860 3519
rect 14948 3283 15184 3519
rect 15272 3283 15508 3519
rect 15596 3283 15832 3519
rect 15920 3283 16156 3519
rect 16244 3283 16480 3519
rect 16568 3283 16804 3519
rect 16892 3283 17128 3519
rect 17216 3283 17452 3519
rect 17540 3283 17776 3519
rect 17864 3283 18100 3519
rect 18188 3283 18424 3519
rect 18512 3283 18748 3519
rect 14300 2952 14536 3188
rect 14624 2952 14860 3188
rect 14948 2952 15184 3188
rect 15272 2952 15508 3188
rect 15596 2952 15832 3188
rect 15920 2952 16156 3188
rect 16244 2952 16480 3188
rect 16568 2952 16804 3188
rect 16892 2952 17128 3188
rect 17216 2952 17452 3188
rect 17540 2952 17776 3188
rect 17864 2952 18100 3188
rect 18188 2952 18424 3188
rect 18512 2952 18748 3188
rect 14300 2621 14536 2857
rect 14624 2621 14860 2857
rect 14948 2621 15184 2857
rect 15272 2621 15508 2857
rect 15596 2621 15832 2857
rect 15920 2621 16156 2857
rect 16244 2621 16480 2857
rect 16568 2621 16804 2857
rect 16892 2621 17128 2857
rect 17216 2621 17452 2857
rect 17540 2621 17776 2857
rect 17864 2621 18100 2857
rect 18188 2621 18424 2857
rect 18512 2621 18748 2857
rect 14300 2290 14536 2526
rect 14624 2290 14860 2526
rect 14948 2290 15184 2526
rect 15272 2290 15508 2526
rect 15596 2290 15832 2526
rect 15920 2290 16156 2526
rect 16244 2290 16480 2526
rect 16568 2290 16804 2526
rect 16892 2290 17128 2526
rect 17216 2290 17452 2526
rect 17540 2290 17776 2526
rect 17864 2290 18100 2526
rect 18188 2290 18424 2526
rect 18512 2290 18748 2526
rect 14300 1959 14536 2195
rect 14624 1959 14860 2195
rect 14948 1959 15184 2195
rect 15272 1959 15508 2195
rect 15596 1959 15832 2195
rect 15920 1959 16156 2195
rect 16244 1959 16480 2195
rect 16568 1959 16804 2195
rect 16892 1959 17128 2195
rect 17216 1959 17452 2195
rect 17540 1959 17776 2195
rect 17864 1959 18100 2195
rect 18188 1959 18424 2195
rect 18512 1959 18748 2195
rect 14300 1628 14536 1864
rect 14624 1628 14860 1864
rect 14948 1628 15184 1864
rect 15272 1628 15508 1864
rect 15596 1628 15832 1864
rect 15920 1628 16156 1864
rect 16244 1628 16480 1864
rect 16568 1628 16804 1864
rect 16892 1628 17128 1864
rect 17216 1628 17452 1864
rect 17540 1628 17776 1864
rect 17864 1628 18100 1864
rect 18188 1628 18424 1864
rect 18512 1628 18748 1864
rect 14300 1297 14536 1533
rect 14624 1297 14860 1533
rect 14948 1297 15184 1533
rect 15272 1297 15508 1533
rect 15596 1297 15832 1533
rect 15920 1297 16156 1533
rect 16244 1297 16480 1533
rect 16568 1297 16804 1533
rect 16892 1297 17128 1533
rect 17216 1297 17452 1533
rect 17540 1297 17776 1533
rect 17864 1297 18100 1533
rect 18188 1297 18424 1533
rect 18512 1297 18748 1533
rect 14300 966 14536 1202
rect 14624 966 14860 1202
rect 14948 966 15184 1202
rect 15272 966 15508 1202
rect 15596 966 15832 1202
rect 15920 966 16156 1202
rect 16244 966 16480 1202
rect 16568 966 16804 1202
rect 16892 966 17128 1202
rect 17216 966 17452 1202
rect 17540 966 17776 1202
rect 17864 966 18100 1202
rect 18188 966 18424 1202
rect 18512 966 18748 1202
rect 14300 635 14536 871
rect 14624 635 14860 871
rect 14948 635 15184 871
rect 15272 635 15508 871
rect 15596 635 15832 871
rect 15920 635 16156 871
rect 16244 635 16480 871
rect 16568 635 16804 871
rect 16892 635 17128 871
rect 17216 635 17452 871
rect 17540 635 17776 871
rect 17864 635 18100 871
rect 18188 635 18424 871
rect 18512 635 18748 871
rect 14300 304 14536 540
rect 14624 304 14860 540
rect 14948 304 15184 540
rect 15272 304 15508 540
rect 15596 304 15832 540
rect 15920 304 16156 540
rect 16244 304 16480 540
rect 16568 304 16804 540
rect 16892 304 17128 540
rect 17216 304 17452 540
rect 17540 304 17776 540
rect 17864 304 18100 540
rect 18188 304 18424 540
rect 18512 304 18748 540
rect 35250 8226 35486 8462
rect 35584 8226 35820 8462
rect 35918 8226 36154 8462
rect 36252 8226 36488 8462
rect 36586 8226 36822 8462
rect 36920 8226 37156 8462
rect 37254 8226 37490 8462
rect 37588 8226 37824 8462
rect 37922 8226 38158 8462
rect 38256 8226 38492 8462
rect 38590 8226 38826 8462
rect 38924 8226 39160 8462
rect 39258 8226 39494 8462
rect 39592 8226 39828 8462
rect 35250 7904 35486 8140
rect 35584 7904 35820 8140
rect 35918 7904 36154 8140
rect 36252 7904 36488 8140
rect 36586 7904 36822 8140
rect 36920 7904 37156 8140
rect 37254 7904 37490 8140
rect 37588 7904 37824 8140
rect 37922 7904 38158 8140
rect 38256 7904 38492 8140
rect 38590 7904 38826 8140
rect 38924 7904 39160 8140
rect 39258 7904 39494 8140
rect 39592 7904 39828 8140
rect 35250 7582 35486 7818
rect 35584 7582 35820 7818
rect 35918 7582 36154 7818
rect 36252 7582 36488 7818
rect 36586 7582 36822 7818
rect 36920 7582 37156 7818
rect 37254 7582 37490 7818
rect 37588 7582 37824 7818
rect 37922 7582 38158 7818
rect 38256 7582 38492 7818
rect 38590 7582 38826 7818
rect 38924 7582 39160 7818
rect 39258 7582 39494 7818
rect 39592 7582 39828 7818
rect 35250 7260 35486 7496
rect 35584 7260 35820 7496
rect 35918 7260 36154 7496
rect 36252 7260 36488 7496
rect 36586 7260 36822 7496
rect 36920 7260 37156 7496
rect 37254 7260 37490 7496
rect 37588 7260 37824 7496
rect 37922 7260 38158 7496
rect 38256 7260 38492 7496
rect 38590 7260 38826 7496
rect 38924 7260 39160 7496
rect 39258 7260 39494 7496
rect 39592 7260 39828 7496
rect 35250 6938 35486 7174
rect 35584 6938 35820 7174
rect 35918 6938 36154 7174
rect 36252 6938 36488 7174
rect 36586 6938 36822 7174
rect 36920 6938 37156 7174
rect 37254 6938 37490 7174
rect 37588 6938 37824 7174
rect 37922 6938 38158 7174
rect 38256 6938 38492 7174
rect 38590 6938 38826 7174
rect 38924 6938 39160 7174
rect 39258 6938 39494 7174
rect 39592 6938 39828 7174
rect 35250 6616 35486 6852
rect 35584 6616 35820 6852
rect 35918 6616 36154 6852
rect 36252 6616 36488 6852
rect 36586 6616 36822 6852
rect 36920 6616 37156 6852
rect 37254 6616 37490 6852
rect 37588 6616 37824 6852
rect 37922 6616 38158 6852
rect 38256 6616 38492 6852
rect 38590 6616 38826 6852
rect 38924 6616 39160 6852
rect 39258 6616 39494 6852
rect 39592 6616 39828 6852
rect 35250 6294 35486 6530
rect 35584 6294 35820 6530
rect 35918 6294 36154 6530
rect 36252 6294 36488 6530
rect 36586 6294 36822 6530
rect 36920 6294 37156 6530
rect 37254 6294 37490 6530
rect 37588 6294 37824 6530
rect 37922 6294 38158 6530
rect 38256 6294 38492 6530
rect 38590 6294 38826 6530
rect 38924 6294 39160 6530
rect 39258 6294 39494 6530
rect 39592 6294 39828 6530
rect 35250 5972 35486 6208
rect 35584 5972 35820 6208
rect 35918 5972 36154 6208
rect 36252 5972 36488 6208
rect 36586 5972 36822 6208
rect 36920 5972 37156 6208
rect 37254 5972 37490 6208
rect 37588 5972 37824 6208
rect 37922 5972 38158 6208
rect 38256 5972 38492 6208
rect 38590 5972 38826 6208
rect 38924 5972 39160 6208
rect 39258 5972 39494 6208
rect 39592 5972 39828 6208
rect 35250 5650 35486 5886
rect 35584 5650 35820 5886
rect 35918 5650 36154 5886
rect 36252 5650 36488 5886
rect 36586 5650 36822 5886
rect 36920 5650 37156 5886
rect 37254 5650 37490 5886
rect 37588 5650 37824 5886
rect 37922 5650 38158 5886
rect 38256 5650 38492 5886
rect 38590 5650 38826 5886
rect 38924 5650 39160 5886
rect 39258 5650 39494 5886
rect 39592 5650 39828 5886
rect 35250 5328 35486 5564
rect 35584 5328 35820 5564
rect 35918 5328 36154 5564
rect 36252 5328 36488 5564
rect 36586 5328 36822 5564
rect 36920 5328 37156 5564
rect 37254 5328 37490 5564
rect 37588 5328 37824 5564
rect 37922 5328 38158 5564
rect 38256 5328 38492 5564
rect 38590 5328 38826 5564
rect 38924 5328 39160 5564
rect 39258 5328 39494 5564
rect 39592 5328 39828 5564
rect 35250 5006 35486 5242
rect 35584 5006 35820 5242
rect 35918 5006 36154 5242
rect 36252 5006 36488 5242
rect 36586 5006 36822 5242
rect 36920 5006 37156 5242
rect 37254 5006 37490 5242
rect 37588 5006 37824 5242
rect 37922 5006 38158 5242
rect 38256 5006 38492 5242
rect 38590 5006 38826 5242
rect 38924 5006 39160 5242
rect 39258 5006 39494 5242
rect 39592 5006 39828 5242
rect 35250 4684 35486 4920
rect 35584 4684 35820 4920
rect 35918 4684 36154 4920
rect 36252 4684 36488 4920
rect 36586 4684 36822 4920
rect 36920 4684 37156 4920
rect 37254 4684 37490 4920
rect 37588 4684 37824 4920
rect 37922 4684 38158 4920
rect 38256 4684 38492 4920
rect 38590 4684 38826 4920
rect 38924 4684 39160 4920
rect 39258 4684 39494 4920
rect 39592 4684 39828 4920
rect 35250 4362 35486 4598
rect 35584 4362 35820 4598
rect 35918 4362 36154 4598
rect 36252 4362 36488 4598
rect 36586 4362 36822 4598
rect 36920 4362 37156 4598
rect 37254 4362 37490 4598
rect 37588 4362 37824 4598
rect 37922 4362 38158 4598
rect 38256 4362 38492 4598
rect 38590 4362 38826 4598
rect 38924 4362 39160 4598
rect 39258 4362 39494 4598
rect 39592 4362 39828 4598
rect 35250 4040 35486 4276
rect 35584 4040 35820 4276
rect 35918 4040 36154 4276
rect 36252 4040 36488 4276
rect 36586 4040 36822 4276
rect 36920 4040 37156 4276
rect 37254 4040 37490 4276
rect 37588 4040 37824 4276
rect 37922 4040 38158 4276
rect 38256 4040 38492 4276
rect 38590 4040 38826 4276
rect 38924 4040 39160 4276
rect 39258 4040 39494 4276
rect 39592 4040 39828 4276
rect 35250 3718 35486 3954
rect 35584 3718 35820 3954
rect 35918 3718 36154 3954
rect 36252 3718 36488 3954
rect 36586 3718 36822 3954
rect 36920 3718 37156 3954
rect 37254 3718 37490 3954
rect 37588 3718 37824 3954
rect 37922 3718 38158 3954
rect 38256 3718 38492 3954
rect 38590 3718 38826 3954
rect 38924 3718 39160 3954
rect 39258 3718 39494 3954
rect 39592 3718 39828 3954
rect 35250 3396 35486 3632
rect 35584 3396 35820 3632
rect 35918 3396 36154 3632
rect 36252 3396 36488 3632
rect 36586 3396 36822 3632
rect 36920 3396 37156 3632
rect 37254 3396 37490 3632
rect 37588 3396 37824 3632
rect 37922 3396 38158 3632
rect 38256 3396 38492 3632
rect 38590 3396 38826 3632
rect 38924 3396 39160 3632
rect 39258 3396 39494 3632
rect 39592 3396 39828 3632
rect 35250 3074 35486 3310
rect 35584 3074 35820 3310
rect 35918 3074 36154 3310
rect 36252 3074 36488 3310
rect 36586 3074 36822 3310
rect 36920 3074 37156 3310
rect 37254 3074 37490 3310
rect 37588 3074 37824 3310
rect 37922 3074 38158 3310
rect 38256 3074 38492 3310
rect 38590 3074 38826 3310
rect 38924 3074 39160 3310
rect 39258 3074 39494 3310
rect 39592 3074 39828 3310
rect 35250 2751 35486 2987
rect 35584 2751 35820 2987
rect 35918 2751 36154 2987
rect 36252 2751 36488 2987
rect 36586 2751 36822 2987
rect 36920 2751 37156 2987
rect 37254 2751 37490 2987
rect 37588 2751 37824 2987
rect 37922 2751 38158 2987
rect 38256 2751 38492 2987
rect 38590 2751 38826 2987
rect 38924 2751 39160 2987
rect 39258 2751 39494 2987
rect 39592 2751 39828 2987
rect 35250 2428 35486 2664
rect 35584 2428 35820 2664
rect 35918 2428 36154 2664
rect 36252 2428 36488 2664
rect 36586 2428 36822 2664
rect 36920 2428 37156 2664
rect 37254 2428 37490 2664
rect 37588 2428 37824 2664
rect 37922 2428 38158 2664
rect 38256 2428 38492 2664
rect 38590 2428 38826 2664
rect 38924 2428 39160 2664
rect 39258 2428 39494 2664
rect 39592 2428 39828 2664
rect 35250 2105 35486 2341
rect 35584 2105 35820 2341
rect 35918 2105 36154 2341
rect 36252 2105 36488 2341
rect 36586 2105 36822 2341
rect 36920 2105 37156 2341
rect 37254 2105 37490 2341
rect 37588 2105 37824 2341
rect 37922 2105 38158 2341
rect 38256 2105 38492 2341
rect 38590 2105 38826 2341
rect 38924 2105 39160 2341
rect 39258 2105 39494 2341
rect 39592 2105 39828 2341
rect 35250 1782 35486 2018
rect 35584 1782 35820 2018
rect 35918 1782 36154 2018
rect 36252 1782 36488 2018
rect 36586 1782 36822 2018
rect 36920 1782 37156 2018
rect 37254 1782 37490 2018
rect 37588 1782 37824 2018
rect 37922 1782 38158 2018
rect 38256 1782 38492 2018
rect 38590 1782 38826 2018
rect 38924 1782 39160 2018
rect 39258 1782 39494 2018
rect 39592 1782 39828 2018
rect 35250 1459 35486 1695
rect 35584 1459 35820 1695
rect 35918 1459 36154 1695
rect 36252 1459 36488 1695
rect 36586 1459 36822 1695
rect 36920 1459 37156 1695
rect 37254 1459 37490 1695
rect 37588 1459 37824 1695
rect 37922 1459 38158 1695
rect 38256 1459 38492 1695
rect 38590 1459 38826 1695
rect 38924 1459 39160 1695
rect 39258 1459 39494 1695
rect 39592 1459 39828 1695
rect 35250 1136 35486 1372
rect 35584 1136 35820 1372
rect 35918 1136 36154 1372
rect 36252 1136 36488 1372
rect 36586 1136 36822 1372
rect 36920 1136 37156 1372
rect 37254 1136 37490 1372
rect 37588 1136 37824 1372
rect 37922 1136 38158 1372
rect 38256 1136 38492 1372
rect 38590 1136 38826 1372
rect 38924 1136 39160 1372
rect 39258 1136 39494 1372
rect 39592 1136 39828 1372
rect 35250 813 35486 1049
rect 35584 813 35820 1049
rect 35918 813 36154 1049
rect 36252 813 36488 1049
rect 36586 813 36822 1049
rect 36920 813 37156 1049
rect 37254 813 37490 1049
rect 37588 813 37824 1049
rect 37922 813 38158 1049
rect 38256 813 38492 1049
rect 38590 813 38826 1049
rect 38924 813 39160 1049
rect 39258 813 39494 1049
rect 39592 813 39828 1049
rect 35250 490 35486 726
rect 35584 490 35820 726
rect 35918 490 36154 726
rect 36252 490 36488 726
rect 36586 490 36822 726
rect 36920 490 37156 726
rect 37254 490 37490 726
rect 37588 490 37824 726
rect 37922 490 38158 726
rect 38256 490 38492 726
rect 38590 490 38826 726
rect 38924 490 39160 726
rect 39258 490 39494 726
rect 39592 490 39828 726
rect 35250 167 35486 403
rect 35584 167 35820 403
rect 35918 167 36154 403
rect 36252 167 36488 403
rect 36586 167 36822 403
rect 36920 167 37156 403
rect 37254 167 37490 403
rect 37588 167 37824 403
rect 37922 167 38158 403
rect 38256 167 38492 403
rect 38590 167 38826 403
rect 38924 167 39160 403
rect 39258 167 39494 403
rect 39592 167 39828 403
<< metal5 >>
rect 0 40559 25423 40733
rect 0 40323 287 40559
rect 523 40323 610 40559
rect 846 40323 933 40559
rect 1169 40323 1256 40559
rect 1492 40323 1579 40559
rect 1815 40323 1902 40559
rect 2138 40323 2225 40559
rect 2461 40323 2548 40559
rect 2784 40323 2871 40559
rect 3107 40323 3194 40559
rect 3430 40323 3517 40559
rect 3753 40323 3840 40559
rect 4076 40323 4163 40559
rect 4399 40323 4486 40559
rect 4722 40323 4809 40559
rect 5045 40323 5132 40559
rect 5368 40323 5455 40559
rect 5691 40323 5778 40559
rect 6014 40323 6101 40559
rect 6337 40323 6424 40559
rect 6660 40323 6747 40559
rect 6983 40323 7070 40559
rect 7306 40323 7393 40559
rect 7629 40323 7716 40559
rect 7952 40323 8039 40559
rect 8275 40323 8362 40559
rect 8598 40323 8685 40559
rect 8921 40323 9008 40559
rect 9244 40323 9331 40559
rect 9567 40323 9654 40559
rect 9890 40323 9977 40559
rect 10213 40323 10300 40559
rect 10536 40323 10623 40559
rect 10859 40323 10946 40559
rect 11182 40323 11269 40559
rect 11505 40323 11592 40559
rect 11828 40323 11915 40559
rect 12151 40323 12238 40559
rect 12474 40323 12561 40559
rect 12797 40323 12884 40559
rect 13120 40323 13207 40559
rect 13443 40323 13530 40559
rect 13766 40323 13853 40559
rect 14089 40323 14176 40559
rect 14412 40323 14499 40559
rect 14735 40323 14822 40559
rect 15058 40323 15145 40559
rect 15381 40323 15468 40559
rect 15704 40323 15791 40559
rect 16027 40323 16114 40559
rect 16350 40323 16437 40559
rect 16673 40323 16760 40559
rect 16996 40323 17082 40559
rect 17318 40323 17404 40559
rect 17640 40323 17726 40559
rect 17962 40323 18048 40559
rect 18284 40323 18370 40559
rect 18606 40323 18692 40559
rect 18928 40323 19014 40559
rect 19250 40323 19336 40559
rect 19572 40323 19658 40559
rect 19894 40323 19980 40559
rect 20216 40323 20302 40559
rect 20538 40323 20624 40559
rect 20860 40323 20946 40559
rect 21182 40323 21268 40559
rect 21504 40323 21590 40559
rect 21826 40323 21912 40559
rect 22148 40323 22234 40559
rect 22470 40323 22556 40559
rect 22792 40323 22878 40559
rect 23114 40323 23200 40559
rect 23436 40323 23522 40559
rect 23758 40323 23844 40559
rect 24080 40323 24166 40559
rect 24402 40323 24488 40559
rect 24724 40323 24810 40559
rect 25046 40323 25132 40559
rect 25368 40323 25423 40559
rect 0 40221 25423 40323
rect 0 39985 287 40221
rect 523 39985 610 40221
rect 846 39985 933 40221
rect 1169 39985 1256 40221
rect 1492 39985 1579 40221
rect 1815 39985 1902 40221
rect 2138 39985 2225 40221
rect 2461 39985 2548 40221
rect 2784 39985 2871 40221
rect 3107 39985 3194 40221
rect 3430 39985 3517 40221
rect 3753 39985 3840 40221
rect 4076 39985 4163 40221
rect 4399 39985 4486 40221
rect 4722 39985 4809 40221
rect 5045 39985 5132 40221
rect 5368 39985 5455 40221
rect 5691 39985 5778 40221
rect 6014 39985 6101 40221
rect 6337 39985 6424 40221
rect 6660 39985 6747 40221
rect 6983 39985 7070 40221
rect 7306 39985 7393 40221
rect 7629 39985 7716 40221
rect 7952 39985 8039 40221
rect 8275 39985 8362 40221
rect 8598 39985 8685 40221
rect 8921 39985 9008 40221
rect 9244 39985 9331 40221
rect 9567 39985 9654 40221
rect 9890 39985 9977 40221
rect 10213 39985 10300 40221
rect 10536 39985 10623 40221
rect 10859 39985 10946 40221
rect 11182 39985 11269 40221
rect 11505 39985 11592 40221
rect 11828 39985 11915 40221
rect 12151 39985 12238 40221
rect 12474 39985 12561 40221
rect 12797 39985 12884 40221
rect 13120 39985 13207 40221
rect 13443 39985 13530 40221
rect 13766 39985 13853 40221
rect 14089 39985 14176 40221
rect 14412 39985 14499 40221
rect 14735 39985 14822 40221
rect 15058 39985 15145 40221
rect 15381 39985 15468 40221
rect 15704 39985 15791 40221
rect 16027 39985 16114 40221
rect 16350 39985 16437 40221
rect 16673 39985 16760 40221
rect 16996 39985 17082 40221
rect 17318 39985 17404 40221
rect 17640 39985 17726 40221
rect 17962 39985 18048 40221
rect 18284 39985 18370 40221
rect 18606 39985 18692 40221
rect 18928 39985 19014 40221
rect 19250 39985 19336 40221
rect 19572 39985 19658 40221
rect 19894 39985 19980 40221
rect 20216 39985 20302 40221
rect 20538 39985 20624 40221
rect 20860 39985 20946 40221
rect 21182 39985 21268 40221
rect 21504 39985 21590 40221
rect 21826 39985 21912 40221
rect 22148 39985 22234 40221
rect 22470 39985 22556 40221
rect 22792 39985 22878 40221
rect 23114 39985 23200 40221
rect 23436 39985 23522 40221
rect 23758 39985 23844 40221
rect 24080 39985 24166 40221
rect 24402 39985 24488 40221
rect 24724 39985 24810 40221
rect 25046 39985 25132 40221
rect 25368 39985 25423 40221
rect 0 39924 25423 39985
tri 25423 39924 26232 40733 sw
rect 0 39900 26232 39924
rect 0 39883 25792 39900
rect 0 39647 287 39883
rect 523 39647 610 39883
rect 846 39647 933 39883
rect 1169 39647 1256 39883
rect 1492 39647 1579 39883
rect 1815 39647 1902 39883
rect 2138 39647 2225 39883
rect 2461 39647 2548 39883
rect 2784 39647 2871 39883
rect 3107 39647 3194 39883
rect 3430 39647 3517 39883
rect 3753 39647 3840 39883
rect 4076 39647 4163 39883
rect 4399 39647 4486 39883
rect 4722 39647 4809 39883
rect 5045 39647 5132 39883
rect 5368 39647 5455 39883
rect 5691 39647 5778 39883
rect 6014 39647 6101 39883
rect 6337 39647 6424 39883
rect 6660 39647 6747 39883
rect 6983 39647 7070 39883
rect 7306 39647 7393 39883
rect 7629 39647 7716 39883
rect 7952 39647 8039 39883
rect 8275 39647 8362 39883
rect 8598 39647 8685 39883
rect 8921 39647 9008 39883
rect 9244 39647 9331 39883
rect 9567 39647 9654 39883
rect 9890 39647 9977 39883
rect 10213 39647 10300 39883
rect 10536 39647 10623 39883
rect 10859 39647 10946 39883
rect 11182 39647 11269 39883
rect 11505 39647 11592 39883
rect 11828 39647 11915 39883
rect 12151 39647 12238 39883
rect 12474 39647 12561 39883
rect 12797 39647 12884 39883
rect 13120 39647 13207 39883
rect 13443 39647 13530 39883
rect 13766 39647 13853 39883
rect 14089 39647 14176 39883
rect 14412 39647 14499 39883
rect 14735 39647 14822 39883
rect 15058 39647 15145 39883
rect 15381 39647 15468 39883
rect 15704 39647 15791 39883
rect 16027 39647 16114 39883
rect 16350 39647 16437 39883
rect 16673 39647 16760 39883
rect 16996 39647 17082 39883
rect 17318 39647 17404 39883
rect 17640 39647 17726 39883
rect 17962 39647 18048 39883
rect 18284 39647 18370 39883
rect 18606 39647 18692 39883
rect 18928 39647 19014 39883
rect 19250 39647 19336 39883
rect 19572 39647 19658 39883
rect 19894 39647 19980 39883
rect 20216 39647 20302 39883
rect 20538 39647 20624 39883
rect 20860 39647 20946 39883
rect 21182 39647 21268 39883
rect 21504 39647 21590 39883
rect 21826 39647 21912 39883
rect 22148 39647 22234 39883
rect 22470 39647 22556 39883
rect 22792 39647 22878 39883
rect 23114 39647 23200 39883
rect 23436 39647 23522 39883
rect 23758 39647 23844 39883
rect 24080 39647 24166 39883
rect 24402 39647 24488 39883
rect 24724 39647 24810 39883
rect 25046 39647 25132 39883
rect 25368 39664 25792 39883
rect 26028 39664 26232 39900
rect 25368 39647 26232 39664
rect 0 39564 26232 39647
rect 0 39545 25792 39564
rect 0 39309 287 39545
rect 523 39309 610 39545
rect 846 39309 933 39545
rect 1169 39309 1256 39545
rect 1492 39309 1579 39545
rect 1815 39309 1902 39545
rect 2138 39309 2225 39545
rect 2461 39309 2548 39545
rect 2784 39309 2871 39545
rect 3107 39309 3194 39545
rect 3430 39309 3517 39545
rect 3753 39309 3840 39545
rect 4076 39309 4163 39545
rect 4399 39309 4486 39545
rect 4722 39309 4809 39545
rect 5045 39309 5132 39545
rect 5368 39309 5455 39545
rect 5691 39309 5778 39545
rect 6014 39309 6101 39545
rect 6337 39309 6424 39545
rect 6660 39309 6747 39545
rect 6983 39309 7070 39545
rect 7306 39309 7393 39545
rect 7629 39309 7716 39545
rect 7952 39309 8039 39545
rect 8275 39309 8362 39545
rect 8598 39309 8685 39545
rect 8921 39309 9008 39545
rect 9244 39309 9331 39545
rect 9567 39309 9654 39545
rect 9890 39309 9977 39545
rect 10213 39309 10300 39545
rect 10536 39309 10623 39545
rect 10859 39309 10946 39545
rect 11182 39309 11269 39545
rect 11505 39309 11592 39545
rect 11828 39309 11915 39545
rect 12151 39309 12238 39545
rect 12474 39309 12561 39545
rect 12797 39309 12884 39545
rect 13120 39309 13207 39545
rect 13443 39309 13530 39545
rect 13766 39309 13853 39545
rect 14089 39309 14176 39545
rect 14412 39309 14499 39545
rect 14735 39309 14822 39545
rect 15058 39309 15145 39545
rect 15381 39309 15468 39545
rect 15704 39309 15791 39545
rect 16027 39309 16114 39545
rect 16350 39309 16437 39545
rect 16673 39309 16760 39545
rect 16996 39309 17082 39545
rect 17318 39309 17404 39545
rect 17640 39309 17726 39545
rect 17962 39309 18048 39545
rect 18284 39309 18370 39545
rect 18606 39309 18692 39545
rect 18928 39309 19014 39545
rect 19250 39309 19336 39545
rect 19572 39309 19658 39545
rect 19894 39309 19980 39545
rect 20216 39309 20302 39545
rect 20538 39309 20624 39545
rect 20860 39309 20946 39545
rect 21182 39309 21268 39545
rect 21504 39309 21590 39545
rect 21826 39309 21912 39545
rect 22148 39309 22234 39545
rect 22470 39309 22556 39545
rect 22792 39309 22878 39545
rect 23114 39309 23200 39545
rect 23436 39309 23522 39545
rect 23758 39309 23844 39545
rect 24080 39309 24166 39545
rect 24402 39309 24488 39545
rect 24724 39309 24810 39545
rect 25046 39309 25132 39545
rect 25368 39328 25792 39545
rect 26028 39328 26232 39564
rect 25368 39309 26232 39328
rect 0 39228 26232 39309
rect 0 39207 25792 39228
rect 0 38971 287 39207
rect 523 38971 610 39207
rect 846 38971 933 39207
rect 1169 38971 1256 39207
rect 1492 38971 1579 39207
rect 1815 38971 1902 39207
rect 2138 38971 2225 39207
rect 2461 38971 2548 39207
rect 2784 38971 2871 39207
rect 3107 38971 3194 39207
rect 3430 38971 3517 39207
rect 3753 38971 3840 39207
rect 4076 38971 4163 39207
rect 4399 38971 4486 39207
rect 4722 38971 4809 39207
rect 5045 38971 5132 39207
rect 5368 38971 5455 39207
rect 5691 38971 5778 39207
rect 6014 38971 6101 39207
rect 6337 38971 6424 39207
rect 6660 38971 6747 39207
rect 6983 38971 7070 39207
rect 7306 38971 7393 39207
rect 7629 38971 7716 39207
rect 7952 38971 8039 39207
rect 8275 38971 8362 39207
rect 8598 38971 8685 39207
rect 8921 38971 9008 39207
rect 9244 38971 9331 39207
rect 9567 38971 9654 39207
rect 9890 38971 9977 39207
rect 10213 38971 10300 39207
rect 10536 38971 10623 39207
rect 10859 38971 10946 39207
rect 11182 38971 11269 39207
rect 11505 38971 11592 39207
rect 11828 38971 11915 39207
rect 12151 38971 12238 39207
rect 12474 38971 12561 39207
rect 12797 38971 12884 39207
rect 13120 38971 13207 39207
rect 13443 38971 13530 39207
rect 13766 38971 13853 39207
rect 14089 38971 14176 39207
rect 14412 38971 14499 39207
rect 14735 38971 14822 39207
rect 15058 38971 15145 39207
rect 15381 38971 15468 39207
rect 15704 38971 15791 39207
rect 16027 38971 16114 39207
rect 16350 38971 16437 39207
rect 16673 38971 16760 39207
rect 16996 38971 17082 39207
rect 17318 38971 17404 39207
rect 17640 38971 17726 39207
rect 17962 38971 18048 39207
rect 18284 38971 18370 39207
rect 18606 38971 18692 39207
rect 18928 38971 19014 39207
rect 19250 38971 19336 39207
rect 19572 38971 19658 39207
rect 19894 38971 19980 39207
rect 20216 38971 20302 39207
rect 20538 38971 20624 39207
rect 20860 38971 20946 39207
rect 21182 38971 21268 39207
rect 21504 38971 21590 39207
rect 21826 38971 21912 39207
rect 22148 38971 22234 39207
rect 22470 38971 22556 39207
rect 22792 38971 22878 39207
rect 23114 38971 23200 39207
rect 23436 38971 23522 39207
rect 23758 38971 23844 39207
rect 24080 38971 24166 39207
rect 24402 38971 24488 39207
rect 24724 38971 24810 39207
rect 25046 38971 25132 39207
rect 25368 38992 25792 39207
rect 26028 38992 26232 39228
rect 25368 38985 26232 38992
tri 26232 38985 27171 39924 sw
rect 25368 38971 27171 38985
rect 0 38961 27171 38971
rect 0 38892 26637 38961
rect 0 38869 25792 38892
rect 0 38633 287 38869
rect 523 38633 610 38869
rect 846 38633 933 38869
rect 1169 38633 1256 38869
rect 1492 38633 1579 38869
rect 1815 38633 1902 38869
rect 2138 38633 2225 38869
rect 2461 38633 2548 38869
rect 2784 38633 2871 38869
rect 3107 38633 3194 38869
rect 3430 38633 3517 38869
rect 3753 38633 3840 38869
rect 4076 38633 4163 38869
rect 4399 38633 4486 38869
rect 4722 38633 4809 38869
rect 5045 38633 5132 38869
rect 5368 38633 5455 38869
rect 5691 38633 5778 38869
rect 6014 38633 6101 38869
rect 6337 38633 6424 38869
rect 6660 38633 6747 38869
rect 6983 38633 7070 38869
rect 7306 38633 7393 38869
rect 7629 38633 7716 38869
rect 7952 38633 8039 38869
rect 8275 38633 8362 38869
rect 8598 38633 8685 38869
rect 8921 38633 9008 38869
rect 9244 38633 9331 38869
rect 9567 38633 9654 38869
rect 9890 38633 9977 38869
rect 10213 38633 10300 38869
rect 10536 38633 10623 38869
rect 10859 38633 10946 38869
rect 11182 38633 11269 38869
rect 11505 38633 11592 38869
rect 11828 38633 11915 38869
rect 12151 38633 12238 38869
rect 12474 38633 12561 38869
rect 12797 38633 12884 38869
rect 13120 38633 13207 38869
rect 13443 38633 13530 38869
rect 13766 38633 13853 38869
rect 14089 38633 14176 38869
rect 14412 38633 14499 38869
rect 14735 38633 14822 38869
rect 15058 38633 15145 38869
rect 15381 38633 15468 38869
rect 15704 38633 15791 38869
rect 16027 38633 16114 38869
rect 16350 38633 16437 38869
rect 16673 38633 16760 38869
rect 16996 38633 17082 38869
rect 17318 38633 17404 38869
rect 17640 38633 17726 38869
rect 17962 38633 18048 38869
rect 18284 38633 18370 38869
rect 18606 38633 18692 38869
rect 18928 38633 19014 38869
rect 19250 38633 19336 38869
rect 19572 38633 19658 38869
rect 19894 38633 19980 38869
rect 20216 38633 20302 38869
rect 20538 38633 20624 38869
rect 20860 38633 20946 38869
rect 21182 38633 21268 38869
rect 21504 38633 21590 38869
rect 21826 38633 21912 38869
rect 22148 38633 22234 38869
rect 22470 38633 22556 38869
rect 22792 38633 22878 38869
rect 23114 38633 23200 38869
rect 23436 38633 23522 38869
rect 23758 38633 23844 38869
rect 24080 38633 24166 38869
rect 24402 38633 24488 38869
rect 24724 38633 24810 38869
rect 25046 38633 25132 38869
rect 25368 38656 25792 38869
rect 26028 38725 26637 38892
rect 26873 38725 27171 38961
rect 26028 38656 27171 38725
rect 25368 38633 27171 38656
rect 0 38625 27171 38633
rect 0 38556 26637 38625
rect 0 38531 25792 38556
rect 0 38295 287 38531
rect 523 38295 610 38531
rect 846 38295 933 38531
rect 1169 38295 1256 38531
rect 1492 38295 1579 38531
rect 1815 38295 1902 38531
rect 2138 38295 2225 38531
rect 2461 38295 2548 38531
rect 2784 38295 2871 38531
rect 3107 38295 3194 38531
rect 3430 38295 3517 38531
rect 3753 38295 3840 38531
rect 4076 38295 4163 38531
rect 4399 38295 4486 38531
rect 4722 38295 4809 38531
rect 5045 38295 5132 38531
rect 5368 38295 5455 38531
rect 5691 38295 5778 38531
rect 6014 38295 6101 38531
rect 6337 38295 6424 38531
rect 6660 38295 6747 38531
rect 6983 38295 7070 38531
rect 7306 38295 7393 38531
rect 7629 38295 7716 38531
rect 7952 38295 8039 38531
rect 8275 38295 8362 38531
rect 8598 38295 8685 38531
rect 8921 38295 9008 38531
rect 9244 38295 9331 38531
rect 9567 38295 9654 38531
rect 9890 38295 9977 38531
rect 10213 38295 10300 38531
rect 10536 38295 10623 38531
rect 10859 38295 10946 38531
rect 11182 38295 11269 38531
rect 11505 38295 11592 38531
rect 11828 38295 11915 38531
rect 12151 38295 12238 38531
rect 12474 38295 12561 38531
rect 12797 38295 12884 38531
rect 13120 38295 13207 38531
rect 13443 38295 13530 38531
rect 13766 38295 13853 38531
rect 14089 38295 14176 38531
rect 14412 38295 14499 38531
rect 14735 38295 14822 38531
rect 15058 38295 15145 38531
rect 15381 38295 15468 38531
rect 15704 38295 15791 38531
rect 16027 38295 16114 38531
rect 16350 38295 16437 38531
rect 16673 38295 16760 38531
rect 16996 38295 17082 38531
rect 17318 38295 17404 38531
rect 17640 38295 17726 38531
rect 17962 38295 18048 38531
rect 18284 38295 18370 38531
rect 18606 38295 18692 38531
rect 18928 38295 19014 38531
rect 19250 38295 19336 38531
rect 19572 38295 19658 38531
rect 19894 38295 19980 38531
rect 20216 38295 20302 38531
rect 20538 38295 20624 38531
rect 20860 38295 20946 38531
rect 21182 38295 21268 38531
rect 21504 38295 21590 38531
rect 21826 38295 21912 38531
rect 22148 38295 22234 38531
rect 22470 38295 22556 38531
rect 22792 38295 22878 38531
rect 23114 38295 23200 38531
rect 23436 38295 23522 38531
rect 23758 38295 23844 38531
rect 24080 38295 24166 38531
rect 24402 38295 24488 38531
rect 24724 38295 24810 38531
rect 25046 38295 25132 38531
rect 25368 38320 25792 38531
rect 26028 38389 26637 38556
rect 26873 38389 27171 38625
rect 26028 38323 27171 38389
tri 27171 38323 27833 38985 sw
rect 26028 38320 27833 38323
rect 25368 38299 27833 38320
rect 25368 38295 27393 38299
rect 0 38289 27393 38295
rect 0 38220 26637 38289
rect 0 38193 25792 38220
rect 0 37957 287 38193
rect 523 37957 610 38193
rect 846 37957 933 38193
rect 1169 37957 1256 38193
rect 1492 37957 1579 38193
rect 1815 37957 1902 38193
rect 2138 37957 2225 38193
rect 2461 37957 2548 38193
rect 2784 37957 2871 38193
rect 3107 37957 3194 38193
rect 3430 37957 3517 38193
rect 3753 37957 3840 38193
rect 4076 37957 4163 38193
rect 4399 37957 4486 38193
rect 4722 37957 4809 38193
rect 5045 37957 5132 38193
rect 5368 37957 5455 38193
rect 5691 37957 5778 38193
rect 6014 37957 6101 38193
rect 6337 37957 6424 38193
rect 6660 37957 6747 38193
rect 6983 37957 7070 38193
rect 7306 37957 7393 38193
rect 7629 37957 7716 38193
rect 7952 37957 8039 38193
rect 8275 37957 8362 38193
rect 8598 37957 8685 38193
rect 8921 37957 9008 38193
rect 9244 37957 9331 38193
rect 9567 37957 9654 38193
rect 9890 37957 9977 38193
rect 10213 37957 10300 38193
rect 10536 37957 10623 38193
rect 10859 37957 10946 38193
rect 11182 37957 11269 38193
rect 11505 37957 11592 38193
rect 11828 37957 11915 38193
rect 12151 37957 12238 38193
rect 12474 37957 12561 38193
rect 12797 37957 12884 38193
rect 13120 37957 13207 38193
rect 13443 37957 13530 38193
rect 13766 37957 13853 38193
rect 14089 37957 14176 38193
rect 14412 37957 14499 38193
rect 14735 37957 14822 38193
rect 15058 37957 15145 38193
rect 15381 37957 15468 38193
rect 15704 37957 15791 38193
rect 16027 37957 16114 38193
rect 16350 37957 16437 38193
rect 16673 37957 16760 38193
rect 16996 37957 17082 38193
rect 17318 37957 17404 38193
rect 17640 37957 17726 38193
rect 17962 37957 18048 38193
rect 18284 37957 18370 38193
rect 18606 37957 18692 38193
rect 18928 37957 19014 38193
rect 19250 37957 19336 38193
rect 19572 37957 19658 38193
rect 19894 37957 19980 38193
rect 20216 37957 20302 38193
rect 20538 37957 20624 38193
rect 20860 37957 20946 38193
rect 21182 37957 21268 38193
rect 21504 37957 21590 38193
rect 21826 37957 21912 38193
rect 22148 37957 22234 38193
rect 22470 37957 22556 38193
rect 22792 37957 22878 38193
rect 23114 37957 23200 38193
rect 23436 37957 23522 38193
rect 23758 37957 23844 38193
rect 24080 37957 24166 38193
rect 24402 37957 24488 38193
rect 24724 37957 24810 38193
rect 25046 37957 25132 38193
rect 25368 37984 25792 38193
rect 26028 38053 26637 38220
rect 26873 38063 27393 38289
rect 27629 38063 27833 38299
rect 26873 38053 27833 38063
rect 26028 37984 27833 38053
rect 25368 37963 27833 37984
rect 25368 37957 27393 37963
rect 0 37953 27393 37957
rect 0 37884 26637 37953
rect 0 37855 25792 37884
rect 0 37619 287 37855
rect 523 37619 610 37855
rect 846 37619 933 37855
rect 1169 37619 1256 37855
rect 1492 37619 1579 37855
rect 1815 37619 1902 37855
rect 2138 37619 2225 37855
rect 2461 37619 2548 37855
rect 2784 37619 2871 37855
rect 3107 37619 3194 37855
rect 3430 37619 3517 37855
rect 3753 37619 3840 37855
rect 4076 37619 4163 37855
rect 4399 37619 4486 37855
rect 4722 37619 4809 37855
rect 5045 37619 5132 37855
rect 5368 37619 5455 37855
rect 5691 37619 5778 37855
rect 6014 37619 6101 37855
rect 6337 37619 6424 37855
rect 6660 37619 6747 37855
rect 6983 37619 7070 37855
rect 7306 37619 7393 37855
rect 7629 37619 7716 37855
rect 7952 37619 8039 37855
rect 8275 37619 8362 37855
rect 8598 37619 8685 37855
rect 8921 37619 9008 37855
rect 9244 37619 9331 37855
rect 9567 37619 9654 37855
rect 9890 37619 9977 37855
rect 10213 37619 10300 37855
rect 10536 37619 10623 37855
rect 10859 37619 10946 37855
rect 11182 37619 11269 37855
rect 11505 37619 11592 37855
rect 11828 37619 11915 37855
rect 12151 37619 12238 37855
rect 12474 37619 12561 37855
rect 12797 37619 12884 37855
rect 13120 37619 13207 37855
rect 13443 37619 13530 37855
rect 13766 37619 13853 37855
rect 14089 37619 14176 37855
rect 14412 37619 14499 37855
rect 14735 37619 14822 37855
rect 15058 37619 15145 37855
rect 15381 37619 15468 37855
rect 15704 37619 15791 37855
rect 16027 37619 16114 37855
rect 16350 37619 16437 37855
rect 16673 37619 16760 37855
rect 16996 37619 17082 37855
rect 17318 37619 17404 37855
rect 17640 37619 17726 37855
rect 17962 37619 18048 37855
rect 18284 37619 18370 37855
rect 18606 37619 18692 37855
rect 18928 37619 19014 37855
rect 19250 37619 19336 37855
rect 19572 37619 19658 37855
rect 19894 37619 19980 37855
rect 20216 37619 20302 37855
rect 20538 37619 20624 37855
rect 20860 37619 20946 37855
rect 21182 37619 21268 37855
rect 21504 37619 21590 37855
rect 21826 37619 21912 37855
rect 22148 37619 22234 37855
rect 22470 37619 22556 37855
rect 22792 37619 22878 37855
rect 23114 37619 23200 37855
rect 23436 37619 23522 37855
rect 23758 37619 23844 37855
rect 24080 37619 24166 37855
rect 24402 37619 24488 37855
rect 24724 37619 24810 37855
rect 25046 37619 25132 37855
rect 25368 37648 25792 37855
rect 26028 37717 26637 37884
rect 26873 37727 27393 37953
rect 27629 37727 27833 37963
rect 26873 37717 27833 37727
rect 26028 37648 27833 37717
rect 25368 37627 27833 37648
rect 25368 37619 27393 37627
rect 0 37617 27393 37619
rect 0 37548 26637 37617
rect 0 37517 25792 37548
rect 0 37281 287 37517
rect 523 37281 610 37517
rect 846 37281 933 37517
rect 1169 37281 1256 37517
rect 1492 37281 1579 37517
rect 1815 37281 1902 37517
rect 2138 37281 2225 37517
rect 2461 37281 2548 37517
rect 2784 37281 2871 37517
rect 3107 37281 3194 37517
rect 3430 37281 3517 37517
rect 3753 37281 3840 37517
rect 4076 37281 4163 37517
rect 4399 37281 4486 37517
rect 4722 37281 4809 37517
rect 5045 37281 5132 37517
rect 5368 37281 5455 37517
rect 5691 37281 5778 37517
rect 6014 37281 6101 37517
rect 6337 37281 6424 37517
rect 6660 37281 6747 37517
rect 6983 37281 7070 37517
rect 7306 37281 7393 37517
rect 7629 37281 7716 37517
rect 7952 37281 8039 37517
rect 8275 37281 8362 37517
rect 8598 37281 8685 37517
rect 8921 37281 9008 37517
rect 9244 37281 9331 37517
rect 9567 37281 9654 37517
rect 9890 37281 9977 37517
rect 10213 37281 10300 37517
rect 10536 37281 10623 37517
rect 10859 37281 10946 37517
rect 11182 37281 11269 37517
rect 11505 37281 11592 37517
rect 11828 37281 11915 37517
rect 12151 37281 12238 37517
rect 12474 37281 12561 37517
rect 12797 37281 12884 37517
rect 13120 37281 13207 37517
rect 13443 37281 13530 37517
rect 13766 37281 13853 37517
rect 14089 37281 14176 37517
rect 14412 37281 14499 37517
rect 14735 37281 14822 37517
rect 15058 37281 15145 37517
rect 15381 37281 15468 37517
rect 15704 37281 15791 37517
rect 16027 37281 16114 37517
rect 16350 37281 16437 37517
rect 16673 37281 16760 37517
rect 16996 37281 17082 37517
rect 17318 37281 17404 37517
rect 17640 37281 17726 37517
rect 17962 37281 18048 37517
rect 18284 37281 18370 37517
rect 18606 37281 18692 37517
rect 18928 37281 19014 37517
rect 19250 37281 19336 37517
rect 19572 37281 19658 37517
rect 19894 37281 19980 37517
rect 20216 37281 20302 37517
rect 20538 37281 20624 37517
rect 20860 37281 20946 37517
rect 21182 37281 21268 37517
rect 21504 37281 21590 37517
rect 21826 37281 21912 37517
rect 22148 37281 22234 37517
rect 22470 37281 22556 37517
rect 22792 37281 22878 37517
rect 23114 37281 23200 37517
rect 23436 37281 23522 37517
rect 23758 37281 23844 37517
rect 24080 37281 24166 37517
rect 24402 37281 24488 37517
rect 24724 37281 24810 37517
rect 25046 37281 25132 37517
rect 25368 37312 25792 37517
rect 26028 37381 26637 37548
rect 26873 37391 27393 37617
rect 27629 37391 27833 37627
rect 26873 37384 27833 37391
tri 27833 37384 28772 38323 sw
rect 26873 37381 28772 37384
rect 26028 37360 28772 37381
rect 26028 37312 28238 37360
rect 25368 37291 28238 37312
rect 25368 37281 27393 37291
rect 0 37211 26637 37281
rect 0 37179 25792 37211
rect 0 36943 287 37179
rect 523 36943 610 37179
rect 846 36943 933 37179
rect 1169 36943 1256 37179
rect 1492 36943 1579 37179
rect 1815 36943 1902 37179
rect 2138 36943 2225 37179
rect 2461 36943 2548 37179
rect 2784 36943 2871 37179
rect 3107 36943 3194 37179
rect 3430 36943 3517 37179
rect 3753 36943 3840 37179
rect 4076 36943 4163 37179
rect 4399 36943 4486 37179
rect 4722 36943 4809 37179
rect 5045 36943 5132 37179
rect 5368 36943 5455 37179
rect 5691 36943 5778 37179
rect 6014 36943 6101 37179
rect 6337 36943 6424 37179
rect 6660 36943 6747 37179
rect 6983 36943 7070 37179
rect 7306 36943 7393 37179
rect 7629 36943 7716 37179
rect 7952 36943 8039 37179
rect 8275 36943 8362 37179
rect 8598 36943 8685 37179
rect 8921 36943 9008 37179
rect 9244 36943 9331 37179
rect 9567 36943 9654 37179
rect 9890 36943 9977 37179
rect 10213 36943 10300 37179
rect 10536 36943 10623 37179
rect 10859 36943 10946 37179
rect 11182 36943 11269 37179
rect 11505 36943 11592 37179
rect 11828 36943 11915 37179
rect 12151 36943 12238 37179
rect 12474 36943 12561 37179
rect 12797 36943 12884 37179
rect 13120 36943 13207 37179
rect 13443 36943 13530 37179
rect 13766 36943 13853 37179
rect 14089 36943 14176 37179
rect 14412 36943 14499 37179
rect 14735 36943 14822 37179
rect 15058 36943 15145 37179
rect 15381 36943 15468 37179
rect 15704 36943 15791 37179
rect 16027 36943 16114 37179
rect 16350 36943 16437 37179
rect 16673 36943 16760 37179
rect 16996 36943 17082 37179
rect 17318 36943 17404 37179
rect 17640 36943 17726 37179
rect 17962 36943 18048 37179
rect 18284 36943 18370 37179
rect 18606 36943 18692 37179
rect 18928 36943 19014 37179
rect 19250 36943 19336 37179
rect 19572 36943 19658 37179
rect 19894 36943 19980 37179
rect 20216 36943 20302 37179
rect 20538 36943 20624 37179
rect 20860 36943 20946 37179
rect 21182 36943 21268 37179
rect 21504 36943 21590 37179
rect 21826 36943 21912 37179
rect 22148 36943 22234 37179
rect 22470 36943 22556 37179
rect 22792 36943 22878 37179
rect 23114 36943 23200 37179
rect 23436 36943 23522 37179
rect 23758 36943 23844 37179
rect 24080 36943 24166 37179
rect 24402 36943 24488 37179
rect 24724 36943 24810 37179
rect 25046 36943 25132 37179
rect 25368 36975 25792 37179
rect 26028 37045 26637 37211
rect 26873 37055 27393 37281
rect 27629 37124 28238 37291
rect 28474 37124 28772 37360
rect 27629 37055 28772 37124
rect 26873 37045 28772 37055
rect 26028 37024 28772 37045
rect 26028 36975 28238 37024
rect 25368 36955 28238 36975
rect 25368 36945 27393 36955
rect 25368 36943 26637 36945
rect 0 36874 26637 36943
rect 0 36841 25792 36874
rect 0 36605 287 36841
rect 523 36605 610 36841
rect 846 36605 933 36841
rect 1169 36605 1256 36841
rect 1492 36605 1579 36841
rect 1815 36605 1902 36841
rect 2138 36605 2225 36841
rect 2461 36605 2548 36841
rect 2784 36605 2871 36841
rect 3107 36605 3194 36841
rect 3430 36605 3517 36841
rect 3753 36605 3840 36841
rect 4076 36605 4163 36841
rect 4399 36605 4486 36841
rect 4722 36605 4809 36841
rect 5045 36605 5132 36841
rect 5368 36605 5455 36841
rect 5691 36605 5778 36841
rect 6014 36605 6101 36841
rect 6337 36605 6424 36841
rect 6660 36605 6747 36841
rect 6983 36605 7070 36841
rect 7306 36605 7393 36841
rect 7629 36605 7716 36841
rect 7952 36605 8039 36841
rect 8275 36605 8362 36841
rect 8598 36605 8685 36841
rect 8921 36605 9008 36841
rect 9244 36605 9331 36841
rect 9567 36605 9654 36841
rect 9890 36605 9977 36841
rect 10213 36605 10300 36841
rect 10536 36605 10623 36841
rect 10859 36605 10946 36841
rect 11182 36605 11269 36841
rect 11505 36605 11592 36841
rect 11828 36605 11915 36841
rect 12151 36605 12238 36841
rect 12474 36605 12561 36841
rect 12797 36605 12884 36841
rect 13120 36605 13207 36841
rect 13443 36605 13530 36841
rect 13766 36605 13853 36841
rect 14089 36605 14176 36841
rect 14412 36605 14499 36841
rect 14735 36605 14822 36841
rect 15058 36605 15145 36841
rect 15381 36605 15468 36841
rect 15704 36605 15791 36841
rect 16027 36605 16114 36841
rect 16350 36605 16437 36841
rect 16673 36605 16760 36841
rect 16996 36605 17082 36841
rect 17318 36605 17404 36841
rect 17640 36605 17726 36841
rect 17962 36605 18048 36841
rect 18284 36605 18370 36841
rect 18606 36605 18692 36841
rect 18928 36605 19014 36841
rect 19250 36605 19336 36841
rect 19572 36605 19658 36841
rect 19894 36605 19980 36841
rect 20216 36605 20302 36841
rect 20538 36605 20624 36841
rect 20860 36605 20946 36841
rect 21182 36605 21268 36841
rect 21504 36605 21590 36841
rect 21826 36605 21912 36841
rect 22148 36605 22234 36841
rect 22470 36605 22556 36841
rect 22792 36605 22878 36841
rect 23114 36605 23200 36841
rect 23436 36605 23522 36841
rect 23758 36605 23844 36841
rect 24080 36605 24166 36841
rect 24402 36605 24488 36841
rect 24724 36605 24810 36841
rect 25046 36605 25132 36841
rect 25368 36638 25792 36841
rect 26028 36709 26637 36874
rect 26873 36719 27393 36945
rect 27629 36788 28238 36955
rect 28474 36788 28772 37024
rect 27629 36722 28772 36788
tri 28772 36722 29434 37384 sw
rect 27629 36719 29434 36722
rect 26873 36709 29434 36719
rect 26028 36698 29434 36709
rect 26028 36688 28994 36698
rect 26028 36638 28238 36688
rect 25368 36619 28238 36638
rect 25368 36609 27393 36619
rect 25368 36605 26637 36609
rect 0 36537 26637 36605
rect 0 36503 25792 36537
rect 0 36267 287 36503
rect 523 36267 610 36503
rect 846 36267 933 36503
rect 1169 36267 1256 36503
rect 1492 36267 1579 36503
rect 1815 36267 1902 36503
rect 2138 36267 2225 36503
rect 2461 36267 2548 36503
rect 2784 36267 2871 36503
rect 3107 36267 3194 36503
rect 3430 36267 3517 36503
rect 3753 36267 3840 36503
rect 4076 36267 4163 36503
rect 4399 36267 4486 36503
rect 4722 36267 4809 36503
rect 5045 36267 5132 36503
rect 5368 36267 5455 36503
rect 5691 36267 5778 36503
rect 6014 36267 6101 36503
rect 6337 36267 6424 36503
rect 6660 36267 6747 36503
rect 6983 36267 7070 36503
rect 7306 36267 7393 36503
rect 7629 36267 7716 36503
rect 7952 36267 8039 36503
rect 8275 36267 8362 36503
rect 8598 36267 8685 36503
rect 8921 36267 9008 36503
rect 9244 36267 9331 36503
rect 9567 36267 9654 36503
rect 9890 36267 9977 36503
rect 10213 36267 10300 36503
rect 10536 36267 10623 36503
rect 10859 36267 10946 36503
rect 11182 36267 11269 36503
rect 11505 36267 11592 36503
rect 11828 36267 11915 36503
rect 12151 36267 12238 36503
rect 12474 36267 12561 36503
rect 12797 36267 12884 36503
rect 13120 36267 13207 36503
rect 13443 36267 13530 36503
rect 13766 36267 13853 36503
rect 14089 36267 14176 36503
rect 14412 36267 14499 36503
rect 14735 36267 14822 36503
rect 15058 36267 15145 36503
rect 15381 36267 15468 36503
rect 15704 36267 15791 36503
rect 16027 36267 16114 36503
rect 16350 36267 16437 36503
rect 16673 36267 16760 36503
rect 16996 36267 17082 36503
rect 17318 36267 17404 36503
rect 17640 36267 17726 36503
rect 17962 36267 18048 36503
rect 18284 36267 18370 36503
rect 18606 36267 18692 36503
rect 18928 36267 19014 36503
rect 19250 36267 19336 36503
rect 19572 36267 19658 36503
rect 19894 36267 19980 36503
rect 20216 36267 20302 36503
rect 20538 36267 20624 36503
rect 20860 36267 20946 36503
rect 21182 36267 21268 36503
rect 21504 36267 21590 36503
rect 21826 36267 21912 36503
rect 22148 36267 22234 36503
rect 22470 36267 22556 36503
rect 22792 36267 22878 36503
rect 23114 36267 23200 36503
rect 23436 36267 23522 36503
rect 23758 36267 23844 36503
rect 24080 36267 24166 36503
rect 24402 36267 24488 36503
rect 24724 36267 24810 36503
rect 25046 36267 25132 36503
rect 25368 36301 25792 36503
rect 26028 36373 26637 36537
rect 26873 36383 27393 36609
rect 27629 36452 28238 36619
rect 28474 36462 28994 36688
rect 29230 36462 29434 36698
rect 28474 36452 29434 36462
rect 27629 36383 29434 36452
rect 26873 36373 29434 36383
rect 26028 36362 29434 36373
rect 26028 36352 28994 36362
rect 26028 36301 28238 36352
rect 25368 36283 28238 36301
rect 25368 36272 27393 36283
rect 25368 36267 26637 36272
rect 0 36200 26637 36267
rect 0 36165 25792 36200
rect 0 35929 287 36165
rect 523 35929 610 36165
rect 846 35929 933 36165
rect 1169 35929 1256 36165
rect 1492 35929 1579 36165
rect 1815 35929 1902 36165
rect 2138 35929 2225 36165
rect 2461 35929 2548 36165
rect 2784 35929 2871 36165
rect 3107 35929 3194 36165
rect 3430 35929 3517 36165
rect 3753 35929 3840 36165
rect 4076 35929 4163 36165
rect 4399 35929 4486 36165
rect 4722 35929 4809 36165
rect 5045 35929 5132 36165
rect 5368 35929 5455 36165
rect 5691 35929 5778 36165
rect 6014 35929 6101 36165
rect 6337 35929 6424 36165
rect 6660 35929 6747 36165
rect 6983 35929 7070 36165
rect 7306 35929 7393 36165
rect 7629 35929 7716 36165
rect 7952 35929 8039 36165
rect 8275 35929 8362 36165
rect 8598 35929 8685 36165
rect 8921 35929 9008 36165
rect 9244 35929 9331 36165
rect 9567 35929 9654 36165
rect 9890 35929 9977 36165
rect 10213 35929 10300 36165
rect 10536 35929 10623 36165
rect 10859 35929 10946 36165
rect 11182 35929 11269 36165
rect 11505 35929 11592 36165
rect 11828 35929 11915 36165
rect 12151 35929 12238 36165
rect 12474 35929 12561 36165
rect 12797 35929 12884 36165
rect 13120 35929 13207 36165
rect 13443 35929 13530 36165
rect 13766 35929 13853 36165
rect 14089 35929 14176 36165
rect 14412 35929 14499 36165
rect 14735 35929 14822 36165
rect 15058 35929 15145 36165
rect 15381 35929 15468 36165
rect 15704 35929 15791 36165
rect 16027 35929 16114 36165
rect 16350 35929 16437 36165
rect 16673 35929 16760 36165
rect 16996 35929 17082 36165
rect 17318 35929 17404 36165
rect 17640 35929 17726 36165
rect 17962 35929 18048 36165
rect 18284 35929 18370 36165
rect 18606 35929 18692 36165
rect 18928 35929 19014 36165
rect 19250 35929 19336 36165
rect 19572 35929 19658 36165
rect 19894 35929 19980 36165
rect 20216 35929 20302 36165
rect 20538 35929 20624 36165
rect 20860 35929 20946 36165
rect 21182 35929 21268 36165
rect 21504 35929 21590 36165
rect 21826 35929 21912 36165
rect 22148 35929 22234 36165
rect 22470 35929 22556 36165
rect 22792 35929 22878 36165
rect 23114 35929 23200 36165
rect 23436 35929 23522 36165
rect 23758 35929 23844 36165
rect 24080 35929 24166 36165
rect 24402 35929 24488 36165
rect 24724 35929 24810 36165
rect 25046 35929 25132 36165
rect 25368 35964 25792 36165
rect 26028 36036 26637 36200
rect 26873 36047 27393 36272
rect 27629 36116 28238 36283
rect 28474 36126 28994 36352
rect 29230 36126 29434 36362
rect 28474 36116 29434 36126
rect 27629 36047 29434 36116
rect 26873 36036 29434 36047
rect 26028 36026 29434 36036
rect 26028 36016 28994 36026
rect 26028 35964 28238 36016
rect 25368 35947 28238 35964
rect 25368 35935 27393 35947
rect 25368 35929 26637 35935
rect 0 35890 26637 35929
tri 23206 33581 25515 35890 ne
rect 25515 35863 26637 35890
rect 25515 35627 25792 35863
rect 26028 35699 26637 35863
rect 26873 35711 27393 35935
rect 27629 35780 28238 35947
rect 28474 35790 28994 36016
rect 29230 35890 29434 36026
tri 29434 35890 30266 36722 sw
rect 29230 35790 30266 35890
rect 28474 35780 30266 35790
rect 27629 35759 30266 35780
rect 27629 35711 29839 35759
rect 26873 35699 29839 35711
rect 26028 35690 29839 35699
rect 26028 35680 28994 35690
rect 26028 35627 28238 35680
rect 25515 35610 28238 35627
rect 25515 35598 27393 35610
rect 25515 35526 26637 35598
rect 25515 35290 25792 35526
rect 26028 35362 26637 35526
rect 26873 35374 27393 35598
rect 27629 35444 28238 35610
rect 28474 35454 28994 35680
rect 29230 35523 29839 35690
rect 30075 35523 30266 35759
rect 29230 35454 30266 35523
rect 28474 35444 30266 35454
rect 27629 35423 30266 35444
rect 27629 35374 29839 35423
rect 26873 35362 29839 35374
rect 26028 35354 29839 35362
rect 26028 35344 28994 35354
rect 26028 35290 28238 35344
rect 25515 35273 28238 35290
rect 25515 35261 27393 35273
rect 25515 35189 26637 35261
rect 25515 34953 25792 35189
rect 26028 35025 26637 35189
rect 26873 35037 27393 35261
rect 27629 35108 28238 35273
rect 28474 35118 28994 35344
rect 29230 35187 29839 35354
rect 30075 35187 30266 35423
rect 29230 35121 30266 35187
tri 30266 35121 31035 35890 sw
rect 29230 35118 31035 35121
rect 28474 35108 31035 35118
rect 27629 35097 31035 35108
rect 27629 35087 30595 35097
rect 27629 35037 29839 35087
rect 26873 35025 29839 35037
rect 26028 35018 29839 35025
rect 26028 35008 28994 35018
rect 26028 34953 28238 35008
rect 25515 34936 28238 34953
rect 25515 34924 27393 34936
rect 25515 34852 26637 34924
rect 25515 34616 25792 34852
rect 26028 34688 26637 34852
rect 26873 34700 27393 34924
rect 27629 34772 28238 34936
rect 28474 34782 28994 35008
rect 29230 34851 29839 35018
rect 30075 34861 30595 35087
rect 30831 34861 31035 35097
rect 30075 34851 31035 34861
rect 29230 34782 31035 34851
rect 28474 34772 31035 34782
rect 27629 34761 31035 34772
rect 27629 34751 30595 34761
rect 27629 34700 29839 34751
rect 26873 34688 29839 34700
rect 26028 34682 29839 34688
rect 26028 34671 28994 34682
rect 26028 34616 28238 34671
rect 25515 34599 28238 34616
rect 25515 34587 27393 34599
rect 25515 34515 26637 34587
rect 25515 34279 25792 34515
rect 26028 34351 26637 34515
rect 26873 34363 27393 34587
rect 27629 34435 28238 34599
rect 28474 34446 28994 34671
rect 29230 34515 29839 34682
rect 30075 34525 30595 34751
rect 30831 34525 31035 34761
rect 30075 34515 31035 34525
rect 29230 34446 31035 34515
rect 28474 34435 31035 34446
rect 27629 34425 31035 34435
rect 27629 34415 30595 34425
rect 27629 34363 29839 34415
rect 26873 34351 29839 34363
rect 26028 34346 29839 34351
rect 26028 34334 28994 34346
rect 26028 34279 28238 34334
rect 25515 34262 28238 34279
rect 25515 34250 27393 34262
rect 25515 34178 26637 34250
rect 25515 33942 25792 34178
rect 26028 34014 26637 34178
rect 26873 34026 27393 34250
rect 27629 34098 28238 34262
rect 28474 34110 28994 34334
rect 29230 34179 29839 34346
rect 30075 34189 30595 34415
rect 30831 34189 31035 34425
rect 30075 34182 31035 34189
tri 31035 34182 31974 35121 sw
rect 30075 34179 31974 34182
rect 29230 34158 31974 34179
rect 29230 34110 31440 34158
rect 28474 34098 31440 34110
rect 27629 34089 31440 34098
rect 27629 34079 30595 34089
rect 27629 34026 29839 34079
rect 26873 34014 29839 34026
rect 26028 34009 29839 34014
rect 26028 33997 28994 34009
rect 26028 33942 28238 33997
rect 25515 33925 28238 33942
rect 25515 33913 27393 33925
rect 25515 33841 26637 33913
rect 25515 33605 25792 33841
rect 26028 33677 26637 33841
rect 26873 33689 27393 33913
rect 27629 33761 28238 33925
rect 28474 33773 28994 33997
rect 29230 33843 29839 34009
rect 30075 33853 30595 34079
rect 30831 33922 31440 34089
rect 31676 33922 31974 34158
rect 30831 33853 31974 33922
rect 30075 33843 31974 33853
rect 29230 33822 31974 33843
rect 29230 33773 31440 33822
rect 28474 33761 31440 33773
rect 27629 33753 31440 33761
rect 27629 33743 30595 33753
rect 27629 33689 29839 33743
rect 26873 33677 29839 33689
rect 26028 33672 29839 33677
rect 26028 33660 28994 33672
rect 26028 33605 28238 33660
rect 25515 33588 28238 33605
rect 25515 33581 27393 33588
tri 25515 32642 26454 33581 ne
rect 26454 33576 27393 33581
rect 26454 33340 26637 33576
rect 26873 33352 27393 33576
rect 27629 33424 28238 33588
rect 28474 33436 28994 33660
rect 29230 33507 29839 33672
rect 30075 33517 30595 33743
rect 30831 33586 31440 33753
rect 31676 33597 31974 33822
tri 31974 33597 32559 34182 sw
rect 31676 33586 32559 33597
rect 30831 33573 32559 33586
rect 30831 33517 32119 33573
rect 30075 33507 32119 33517
rect 29230 33486 32119 33507
rect 29230 33436 31440 33486
rect 28474 33424 31440 33436
rect 27629 33417 31440 33424
rect 27629 33407 30595 33417
rect 27629 33352 29839 33407
rect 26873 33340 29839 33352
rect 26454 33335 29839 33340
rect 26454 33323 28994 33335
rect 26454 33251 28238 33323
rect 26454 33239 27393 33251
rect 26454 33003 26637 33239
rect 26873 33015 27393 33239
rect 27629 33087 28238 33251
rect 28474 33099 28994 33323
rect 29230 33171 29839 33335
rect 30075 33181 30595 33407
rect 30831 33250 31440 33417
rect 31676 33337 32119 33486
rect 32355 33337 32559 33573
rect 31676 33250 32559 33337
rect 30831 33237 32559 33250
rect 30831 33181 32119 33237
rect 30075 33171 32119 33181
rect 29230 33150 32119 33171
rect 29230 33099 31440 33150
rect 28474 33087 31440 33099
rect 27629 33081 31440 33087
rect 27629 33070 30595 33081
rect 27629 33015 29839 33070
rect 26873 33003 29839 33015
rect 26454 32998 29839 33003
rect 26454 32986 28994 32998
rect 26454 32914 28238 32986
rect 26454 32902 27393 32914
rect 26454 32666 26637 32902
rect 26873 32678 27393 32902
rect 27629 32750 28238 32914
rect 28474 32762 28994 32986
rect 29230 32834 29839 32998
rect 30075 32845 30595 33070
rect 30831 32914 31440 33081
rect 31676 33001 32119 33150
rect 32355 33001 32559 33237
rect 31676 32914 32559 33001
rect 30831 32901 32559 32914
rect 30831 32845 32119 32901
rect 30075 32834 32119 32845
rect 29230 32814 32119 32834
rect 29230 32762 31440 32814
rect 28474 32750 31440 32762
rect 27629 32745 31440 32750
rect 27629 32733 30595 32745
rect 27629 32678 29839 32733
rect 26873 32666 29839 32678
rect 26454 32661 29839 32666
rect 26454 32649 28994 32661
rect 26454 32642 28238 32649
tri 26454 31980 27116 32642 ne
rect 27116 32577 28238 32642
rect 27116 32341 27393 32577
rect 27629 32413 28238 32577
rect 28474 32425 28994 32649
rect 29230 32497 29839 32661
rect 30075 32509 30595 32733
rect 30831 32578 31440 32745
rect 31676 32665 32119 32814
rect 32355 32665 32559 32901
rect 31676 32658 32559 32665
tri 32559 32658 33498 33597 sw
rect 31676 32634 33498 32658
rect 31676 32578 32964 32634
rect 30831 32565 32964 32578
rect 30831 32509 32119 32565
rect 30075 32497 32119 32509
rect 29230 32478 32119 32497
rect 29230 32425 31440 32478
rect 28474 32413 31440 32425
rect 27629 32408 31440 32413
rect 27629 32396 30595 32408
rect 27629 32341 29839 32396
rect 27116 32324 29839 32341
rect 27116 32312 28994 32324
rect 27116 32240 28238 32312
rect 27116 32004 27393 32240
rect 27629 32076 28238 32240
rect 28474 32088 28994 32312
rect 29230 32160 29839 32324
rect 30075 32172 30595 32396
rect 30831 32242 31440 32408
rect 31676 32329 32119 32478
rect 32355 32398 32964 32565
rect 33200 32398 33498 32634
rect 32355 32329 33498 32398
rect 31676 32298 33498 32329
rect 31676 32242 32964 32298
rect 30831 32229 32964 32242
rect 30831 32172 32119 32229
rect 30075 32160 32119 32172
rect 29230 32142 32119 32160
rect 29230 32088 31440 32142
rect 28474 32076 31440 32088
rect 27629 32071 31440 32076
rect 27629 32059 30595 32071
rect 27629 32004 29839 32059
rect 27116 31987 29839 32004
rect 27116 31980 28994 31987
tri 27116 31041 28055 31980 ne
rect 28055 31975 28994 31980
rect 28055 31739 28238 31975
rect 28474 31751 28994 31975
rect 29230 31823 29839 31987
rect 30075 31835 30595 32059
rect 30831 31906 31440 32071
rect 31676 31993 32119 32142
rect 32355 32062 32964 32229
rect 33200 32062 33498 32298
rect 32355 31996 33498 32062
tri 33498 31996 34160 32658 sw
rect 32355 31993 34160 31996
rect 31676 31972 34160 31993
rect 31676 31962 33720 31972
rect 31676 31906 32964 31962
rect 30831 31893 32964 31906
rect 30831 31835 32119 31893
rect 30075 31823 32119 31835
rect 29230 31806 32119 31823
rect 29230 31751 31440 31806
rect 28474 31739 31440 31751
rect 28055 31734 31440 31739
rect 28055 31722 30595 31734
rect 28055 31650 29839 31722
rect 28055 31638 28994 31650
rect 28055 31402 28238 31638
rect 28474 31414 28994 31638
rect 29230 31486 29839 31650
rect 30075 31498 30595 31722
rect 30831 31570 31440 31734
rect 31676 31657 32119 31806
rect 32355 31726 32964 31893
rect 33200 31736 33720 31962
rect 33956 31736 34160 31972
rect 33200 31726 34160 31736
rect 32355 31657 34160 31726
rect 31676 31636 34160 31657
rect 31676 31626 33720 31636
rect 31676 31570 32964 31626
rect 30831 31557 32964 31570
rect 30831 31498 32119 31557
rect 30075 31486 32119 31498
rect 29230 31469 32119 31486
rect 29230 31414 31440 31469
rect 28474 31402 31440 31414
rect 28055 31397 31440 31402
rect 28055 31385 30595 31397
rect 28055 31313 29839 31385
rect 28055 31301 28994 31313
rect 28055 31065 28238 31301
rect 28474 31077 28994 31301
rect 29230 31149 29839 31313
rect 30075 31161 30595 31385
rect 30831 31233 31440 31397
rect 31676 31321 32119 31469
rect 32355 31390 32964 31557
rect 33200 31400 33720 31626
rect 33956 31400 34160 31636
rect 33200 31390 34160 31400
rect 32355 31321 34160 31390
rect 31676 31300 34160 31321
rect 31676 31290 33720 31300
rect 31676 31233 32964 31290
rect 30831 31221 32964 31233
rect 30831 31161 32119 31221
rect 30075 31149 32119 31161
rect 29230 31132 32119 31149
rect 29230 31077 31440 31132
rect 28474 31065 31440 31077
rect 28055 31060 31440 31065
rect 28055 31048 30595 31060
rect 28055 31041 29839 31048
tri 28055 30379 28717 31041 ne
rect 28717 30976 29839 31041
rect 28717 30740 28994 30976
rect 29230 30812 29839 30976
rect 30075 30824 30595 31048
rect 30831 30896 31440 31060
rect 31676 30985 32119 31132
rect 32355 31054 32964 31221
rect 33200 31064 33720 31290
rect 33956 31064 34160 31300
rect 33200 31057 34160 31064
tri 34160 31057 35099 31996 sw
rect 33200 31054 35099 31057
rect 32355 31033 35099 31054
rect 32355 30985 34565 31033
rect 31676 30964 34565 30985
rect 31676 30954 33720 30964
rect 31676 30896 32964 30954
rect 30831 30884 32964 30896
rect 30831 30824 32119 30884
rect 30075 30812 32119 30824
rect 29230 30795 32119 30812
rect 29230 30740 31440 30795
rect 28717 30723 31440 30740
rect 28717 30711 30595 30723
rect 28717 30639 29839 30711
rect 28717 30403 28994 30639
rect 29230 30475 29839 30639
rect 30075 30487 30595 30711
rect 30831 30559 31440 30723
rect 31676 30648 32119 30795
rect 32355 30718 32964 30884
rect 33200 30728 33720 30954
rect 33956 30797 34565 30964
rect 34801 30999 35099 31033
tri 35099 30999 35157 31057 sw
rect 34801 30797 35157 30999
rect 33956 30728 35157 30797
rect 33200 30718 35157 30728
rect 32355 30697 35157 30718
rect 32355 30648 34565 30697
rect 31676 30628 34565 30648
rect 31676 30618 33720 30628
rect 31676 30559 32964 30618
rect 30831 30547 32964 30559
rect 30831 30487 32119 30547
rect 30075 30475 32119 30487
rect 29230 30458 32119 30475
rect 29230 30403 31440 30458
rect 28717 30386 31440 30403
rect 28717 30379 30595 30386
tri 28717 29440 29656 30379 ne
rect 29656 30374 30595 30379
rect 29656 30138 29839 30374
rect 30075 30150 30595 30374
rect 30831 30222 31440 30386
rect 31676 30311 32119 30458
rect 32355 30382 32964 30547
rect 33200 30392 33720 30618
rect 33956 30461 34565 30628
rect 34801 30461 35157 30697
rect 33956 30392 35157 30461
rect 33200 30382 35157 30392
rect 32355 30361 35157 30382
rect 32355 30311 34565 30361
rect 31676 30292 34565 30311
rect 31676 30282 33720 30292
rect 31676 30222 32964 30282
rect 30831 30210 32964 30222
rect 30831 30150 32119 30210
rect 30075 30138 32119 30150
rect 29656 30121 32119 30138
rect 29656 30049 31440 30121
rect 29656 30037 30595 30049
rect 29656 29801 29839 30037
rect 30075 29813 30595 30037
rect 30831 29885 31440 30049
rect 31676 29974 32119 30121
rect 32355 30046 32964 30210
rect 33200 30056 33720 30282
rect 33956 30125 34565 30292
rect 34801 30257 35157 30361
tri 35157 30257 35899 30999 sw
rect 34801 30233 35899 30257
rect 34801 30125 35365 30233
rect 33956 30056 35365 30125
rect 33200 30046 35365 30056
rect 32355 30025 35365 30046
rect 32355 29974 34565 30025
rect 31676 29956 34565 29974
rect 31676 29945 33720 29956
rect 31676 29885 32964 29945
rect 30831 29873 32964 29885
rect 30831 29813 32119 29873
rect 30075 29801 32119 29813
rect 29656 29784 32119 29801
rect 29656 29712 31440 29784
rect 29656 29700 30595 29712
rect 29656 29464 29839 29700
rect 30075 29476 30595 29700
rect 30831 29548 31440 29712
rect 31676 29637 32119 29784
rect 32355 29709 32964 29873
rect 33200 29720 33720 29945
rect 33956 29789 34565 29956
rect 34801 29997 35365 30025
rect 35601 29997 35899 30233
rect 34801 29901 35899 29997
rect 34801 29789 35365 29901
rect 33956 29720 35365 29789
rect 33200 29709 35365 29720
rect 32355 29689 35365 29709
rect 32355 29637 34565 29689
rect 31676 29620 34565 29637
rect 31676 29608 33720 29620
rect 31676 29548 32964 29608
rect 30831 29536 32964 29548
rect 30831 29476 32119 29536
rect 30075 29464 32119 29476
rect 29656 29447 32119 29464
rect 29656 29440 31440 29447
tri 29656 28830 30266 29440 ne
rect 30266 29375 31440 29440
rect 30266 29139 30595 29375
rect 30831 29211 31440 29375
rect 31676 29300 32119 29447
rect 32355 29372 32964 29536
rect 33200 29384 33720 29608
rect 33956 29453 34565 29620
rect 34801 29665 35365 29689
rect 35601 29665 35899 29901
rect 34801 29569 35899 29665
rect 34801 29453 35365 29569
rect 33956 29384 35365 29453
rect 33200 29372 35365 29384
rect 32355 29353 35365 29372
rect 32355 29300 34565 29353
rect 31676 29283 34565 29300
rect 31676 29271 33720 29283
rect 31676 29211 32964 29271
rect 30831 29199 32964 29211
rect 30831 29139 32119 29199
rect 30266 29110 32119 29139
rect 30266 29038 31440 29110
rect 30266 28830 30595 29038
tri 30266 28778 30318 28830 ne
rect 30318 28802 30595 28830
rect 30831 28874 31440 29038
rect 31676 28963 32119 29110
rect 32355 29035 32964 29199
rect 33200 29047 33720 29271
rect 33956 29117 34565 29283
rect 34801 29333 35365 29353
rect 35601 29385 35899 29569
tri 35899 29385 36771 30257 sw
rect 35601 29361 36771 29385
rect 35601 29333 36237 29361
rect 34801 29237 36237 29333
rect 34801 29117 35365 29237
rect 33956 29047 35365 29117
rect 33200 29035 35365 29047
rect 32355 29017 35365 29035
rect 32355 28963 34565 29017
rect 31676 28946 34565 28963
rect 31676 28934 33720 28946
rect 31676 28874 32964 28934
rect 30831 28862 32964 28874
rect 30831 28802 32119 28862
rect 30318 28778 32119 28802
tri 30318 27839 31257 28778 ne
rect 31257 28773 32119 28778
rect 31257 28537 31440 28773
rect 31676 28626 32119 28773
rect 32355 28698 32964 28862
rect 33200 28710 33720 28934
rect 33956 28781 34565 28946
rect 34801 29001 35365 29017
rect 35601 29125 36237 29237
rect 36473 29125 36771 29361
rect 35601 29029 36771 29125
rect 35601 29001 36237 29029
rect 34801 28905 36237 29001
rect 34801 28781 35365 28905
rect 33956 28710 35365 28781
rect 33200 28698 35365 28710
rect 32355 28681 35365 28698
rect 32355 28626 34565 28681
rect 31676 28609 34565 28626
rect 31676 28597 33720 28609
rect 31676 28537 32964 28597
rect 31257 28525 32964 28537
rect 31257 28436 32119 28525
rect 31257 28200 31440 28436
rect 31676 28289 32119 28436
rect 32355 28361 32964 28525
rect 33200 28373 33720 28597
rect 33956 28445 34565 28609
rect 34801 28669 35365 28681
rect 35601 28793 36237 28905
rect 36473 28830 36771 29029
tri 36771 28830 37326 29385 sw
rect 36473 28793 37326 28830
rect 35601 28697 37326 28793
rect 35601 28669 36237 28697
rect 34801 28573 36237 28669
rect 34801 28445 35365 28573
rect 33956 28373 35365 28445
rect 33200 28361 35365 28373
rect 32355 28344 35365 28361
rect 32355 28289 34565 28344
rect 31676 28272 34565 28289
rect 31676 28260 33720 28272
rect 31676 28200 32964 28260
rect 31257 28188 32964 28200
rect 31257 28099 32119 28188
rect 31257 27863 31440 28099
rect 31676 27952 32119 28099
rect 32355 28024 32964 28188
rect 33200 28036 33720 28260
rect 33956 28108 34565 28272
rect 34801 28337 35365 28344
rect 35601 28461 36237 28573
rect 36473 28499 37326 28697
tri 37326 28499 37657 28830 sw
rect 36473 28475 37657 28499
rect 36473 28461 37123 28475
rect 35601 28365 37123 28461
rect 35601 28337 36237 28365
rect 34801 28241 36237 28337
rect 34801 28108 35365 28241
rect 33956 28036 35365 28108
rect 33200 28024 35365 28036
rect 32355 28007 35365 28024
rect 32355 27952 34565 28007
rect 31676 27935 34565 27952
rect 31676 27923 33720 27935
rect 31676 27863 32964 27923
rect 31257 27851 32964 27863
rect 31257 27839 32119 27851
tri 31257 27254 31842 27839 ne
rect 31842 27615 32119 27839
rect 32355 27687 32964 27851
rect 33200 27699 33720 27923
rect 33956 27771 34565 27935
rect 34801 28005 35365 28007
rect 35601 28129 36237 28241
rect 36473 28239 37123 28365
rect 37359 28239 37657 28475
rect 36473 28132 37657 28239
rect 36473 28129 37123 28132
rect 35601 28033 37123 28129
rect 35601 28005 36237 28033
rect 34801 27909 36237 28005
rect 34801 27771 35365 27909
rect 33956 27699 35365 27771
rect 33200 27687 35365 27699
rect 32355 27673 35365 27687
rect 35601 27797 36237 27909
rect 36473 27896 37123 28033
rect 37359 27896 37657 28132
rect 36473 27797 37657 27896
rect 35601 27789 37657 27797
rect 35601 27701 37123 27789
rect 35601 27673 36237 27701
rect 32355 27670 36237 27673
rect 32355 27615 34565 27670
rect 31842 27598 34565 27615
rect 31842 27586 33720 27598
rect 31842 27514 32964 27586
rect 31842 27278 32119 27514
rect 32355 27350 32964 27514
rect 33200 27362 33720 27586
rect 33956 27434 34565 27598
rect 34801 27577 36237 27670
rect 34801 27434 35365 27577
rect 33956 27362 35365 27434
rect 33200 27350 35365 27362
rect 32355 27341 35365 27350
rect 35601 27465 36237 27577
rect 36473 27553 37123 27701
rect 37359 27673 37657 27789
tri 37657 27673 38483 28499 sw
rect 37359 27649 38483 27673
rect 37359 27553 37949 27649
rect 36473 27465 37949 27553
rect 35601 27446 37949 27465
rect 35601 27369 37123 27446
rect 35601 27341 36237 27369
rect 32355 27333 36237 27341
rect 32355 27278 34565 27333
rect 31842 27261 34565 27278
rect 31842 27254 33720 27261
tri 31842 26315 32781 27254 ne
rect 32781 27249 33720 27254
rect 32781 27013 32964 27249
rect 33200 27025 33720 27249
rect 33956 27097 34565 27261
rect 34801 27245 36237 27333
rect 34801 27097 35365 27245
rect 33956 27025 35365 27097
rect 33200 27013 35365 27025
rect 32781 27009 35365 27013
rect 35601 27133 36237 27245
rect 36473 27210 37123 27369
rect 37359 27413 37949 27446
rect 38185 27413 38483 27649
rect 37359 27324 38483 27413
rect 37359 27210 37949 27324
rect 36473 27133 37949 27210
rect 35601 27103 37949 27133
rect 35601 27037 37123 27103
rect 35601 27009 36237 27037
rect 32781 26996 36237 27009
rect 32781 26924 34565 26996
rect 32781 26912 33720 26924
rect 32781 26676 32964 26912
rect 33200 26688 33720 26912
rect 33956 26760 34565 26924
rect 34801 26913 36237 26996
rect 34801 26760 35365 26913
rect 33956 26688 35365 26760
rect 33200 26677 35365 26688
rect 35601 26801 36237 26913
rect 36473 26867 37123 27037
rect 37359 27088 37949 27103
rect 38185 27088 38483 27324
rect 37359 26999 38483 27088
rect 37359 26867 37949 26999
rect 36473 26801 37949 26867
rect 35601 26763 37949 26801
rect 38185 26874 38483 26999
tri 38483 26874 39282 27673 sw
rect 38185 26850 39282 26874
rect 38185 26763 38748 26850
rect 35601 26760 38748 26763
rect 35601 26705 37123 26760
rect 35601 26677 36237 26705
rect 33200 26676 36237 26677
rect 32781 26659 36237 26676
rect 32781 26587 34565 26659
rect 32781 26575 33720 26587
rect 32781 26339 32964 26575
rect 33200 26351 33720 26575
rect 33956 26423 34565 26587
rect 34801 26580 36237 26659
rect 34801 26423 35365 26580
rect 33956 26351 35365 26423
rect 33200 26344 35365 26351
rect 35601 26469 36237 26580
rect 36473 26524 37123 26705
rect 37359 26673 38748 26760
rect 37359 26524 37949 26673
rect 36473 26469 37949 26524
rect 35601 26437 37949 26469
rect 38185 26614 38748 26673
rect 38984 26614 39282 26850
rect 38185 26525 39282 26614
rect 38185 26437 38748 26525
rect 35601 26416 38748 26437
rect 35601 26373 37123 26416
rect 35601 26344 36237 26373
rect 33200 26339 36237 26344
rect 32781 26322 36237 26339
rect 32781 26315 34565 26322
tri 32781 25653 33443 26315 ne
rect 33443 26250 34565 26315
rect 33443 26014 33720 26250
rect 33956 26086 34565 26250
rect 34801 26247 36237 26322
rect 34801 26086 35365 26247
rect 33956 26014 35365 26086
rect 33443 26011 35365 26014
rect 35601 26137 36237 26247
rect 36473 26180 37123 26373
rect 37359 26347 38748 26416
rect 37359 26180 37949 26347
rect 36473 26137 37949 26180
rect 35601 26111 37949 26137
rect 38185 26289 38748 26347
rect 38984 26289 39282 26525
rect 38185 26200 39282 26289
rect 38185 26111 38748 26200
rect 35601 26072 38748 26111
rect 35601 26041 37123 26072
rect 35601 26011 36237 26041
rect 33443 25985 36237 26011
rect 33443 25913 34565 25985
rect 33443 25677 33720 25913
rect 33956 25749 34565 25913
rect 34801 25914 36237 25985
rect 34801 25749 35365 25914
rect 33956 25678 35365 25749
rect 35601 25805 36237 25914
rect 36473 25836 37123 26041
rect 37359 26021 38748 26072
rect 37359 25836 37949 26021
rect 36473 25805 37949 25836
rect 35601 25785 37949 25805
rect 38185 25964 38748 26021
rect 38984 26156 39282 26200
tri 39282 26156 40000 26874 sw
rect 38984 25964 40000 26156
rect 38185 25875 40000 25964
rect 38185 25785 38748 25875
rect 35601 25728 38748 25785
rect 35601 25709 37123 25728
rect 35601 25678 36237 25709
rect 33956 25677 36237 25678
rect 33443 25653 36237 25677
tri 33443 24714 34382 25653 ne
rect 34382 25648 36237 25653
rect 34382 25412 34565 25648
rect 34801 25581 36237 25648
rect 34801 25412 35365 25581
rect 34382 25345 35365 25412
rect 35601 25473 36237 25581
rect 36473 25492 37123 25709
rect 37359 25695 38748 25728
rect 37359 25492 37949 25695
rect 36473 25473 37949 25492
rect 35601 25459 37949 25473
rect 38185 25639 38748 25695
rect 38984 25639 40000 25875
rect 38185 25550 40000 25639
rect 38185 25459 38748 25550
rect 35601 25384 38748 25459
rect 35601 25377 37123 25384
rect 35601 25345 36237 25377
rect 34382 25311 36237 25345
rect 34382 25075 34565 25311
rect 34801 25248 36237 25311
rect 34801 25075 35365 25248
rect 34382 25012 35365 25075
rect 35601 25141 36237 25248
rect 36473 25148 37123 25377
rect 37359 25369 38748 25384
rect 37359 25148 37949 25369
rect 36473 25141 37949 25148
rect 35601 25133 37949 25141
rect 38185 25314 38748 25369
rect 38984 25314 40000 25550
rect 38185 25225 40000 25314
rect 38185 25133 38748 25225
rect 35601 25044 38748 25133
rect 35601 25012 36237 25044
rect 34382 24974 36237 25012
rect 34382 24738 34565 24974
rect 34801 24915 36237 24974
rect 34801 24738 35365 24915
rect 34382 24714 35365 24738
tri 34382 23939 35157 24714 ne
rect 35157 24679 35365 24714
rect 35601 24808 36237 24915
rect 36473 25043 38748 25044
rect 36473 25040 37949 25043
rect 36473 24808 37123 25040
rect 35601 24804 37123 24808
rect 37359 24807 37949 25040
rect 38185 24989 38748 25043
rect 38984 24989 40000 25225
rect 38185 24899 40000 24989
rect 38185 24807 38748 24899
rect 37359 24804 38748 24807
rect 35601 24717 38748 24804
rect 35601 24711 37949 24717
rect 35601 24679 36237 24711
rect 35157 24475 36237 24679
rect 36473 24696 37949 24711
rect 36473 24475 37123 24696
rect 35157 24460 37123 24475
rect 37359 24481 37949 24696
rect 38185 24663 38748 24717
rect 38984 24663 40000 24899
rect 38185 24573 40000 24663
rect 38185 24481 38748 24573
rect 37359 24460 38748 24481
rect 35157 24337 38748 24460
rect 38984 24337 40000 24573
rect 35157 23918 40000 24337
rect 35157 23682 35250 23918
rect 35486 23682 35584 23918
rect 35820 23682 35918 23918
rect 36154 23682 36252 23918
rect 36488 23682 36586 23918
rect 36822 23682 36920 23918
rect 37156 23682 37254 23918
rect 37490 23682 37588 23918
rect 37824 23682 37922 23918
rect 38158 23682 38256 23918
rect 38492 23682 38590 23918
rect 38826 23682 38924 23918
rect 39160 23682 39258 23918
rect 39494 23682 39592 23918
rect 39828 23682 40000 23918
rect 35157 23596 40000 23682
rect 35157 23360 35250 23596
rect 35486 23360 35584 23596
rect 35820 23360 35918 23596
rect 36154 23360 36252 23596
rect 36488 23360 36586 23596
rect 36822 23360 36920 23596
rect 37156 23360 37254 23596
rect 37490 23360 37588 23596
rect 37824 23360 37922 23596
rect 38158 23360 38256 23596
rect 38492 23360 38590 23596
rect 38826 23360 38924 23596
rect 39160 23360 39258 23596
rect 39494 23360 39592 23596
rect 39828 23360 40000 23596
rect 35157 23274 40000 23360
rect 35157 23038 35250 23274
rect 35486 23038 35584 23274
rect 35820 23038 35918 23274
rect 36154 23038 36252 23274
rect 36488 23038 36586 23274
rect 36822 23038 36920 23274
rect 37156 23038 37254 23274
rect 37490 23038 37588 23274
rect 37824 23038 37922 23274
rect 38158 23038 38256 23274
rect 38492 23038 38590 23274
rect 38826 23038 38924 23274
rect 39160 23038 39258 23274
rect 39494 23038 39592 23274
rect 39828 23038 40000 23274
rect 35157 22952 40000 23038
rect 35157 22716 35250 22952
rect 35486 22716 35584 22952
rect 35820 22716 35918 22952
rect 36154 22716 36252 22952
rect 36488 22716 36586 22952
rect 36822 22716 36920 22952
rect 37156 22716 37254 22952
rect 37490 22716 37588 22952
rect 37824 22716 37922 22952
rect 38158 22716 38256 22952
rect 38492 22716 38590 22952
rect 38826 22716 38924 22952
rect 39160 22716 39258 22952
rect 39494 22716 39592 22952
rect 39828 22716 40000 22952
rect 35157 22630 40000 22716
rect 35157 22394 35250 22630
rect 35486 22394 35584 22630
rect 35820 22394 35918 22630
rect 36154 22394 36252 22630
rect 36488 22394 36586 22630
rect 36822 22394 36920 22630
rect 37156 22394 37254 22630
rect 37490 22394 37588 22630
rect 37824 22394 37922 22630
rect 38158 22394 38256 22630
rect 38492 22394 38590 22630
rect 38826 22394 38924 22630
rect 39160 22394 39258 22630
rect 39494 22394 39592 22630
rect 39828 22394 40000 22630
rect 35157 22308 40000 22394
rect 35157 22072 35250 22308
rect 35486 22072 35584 22308
rect 35820 22072 35918 22308
rect 36154 22072 36252 22308
rect 36488 22072 36586 22308
rect 36822 22072 36920 22308
rect 37156 22072 37254 22308
rect 37490 22072 37588 22308
rect 37824 22072 37922 22308
rect 38158 22072 38256 22308
rect 38492 22072 38590 22308
rect 38826 22072 38924 22308
rect 39160 22072 39258 22308
rect 39494 22072 39592 22308
rect 39828 22072 40000 22308
rect 35157 21986 40000 22072
rect 35157 21750 35250 21986
rect 35486 21750 35584 21986
rect 35820 21750 35918 21986
rect 36154 21750 36252 21986
rect 36488 21750 36586 21986
rect 36822 21750 36920 21986
rect 37156 21750 37254 21986
rect 37490 21750 37588 21986
rect 37824 21750 37922 21986
rect 38158 21750 38256 21986
rect 38492 21750 38590 21986
rect 38826 21750 38924 21986
rect 39160 21750 39258 21986
rect 39494 21750 39592 21986
rect 39828 21750 40000 21986
rect 35157 21664 40000 21750
rect 35157 21428 35250 21664
rect 35486 21428 35584 21664
rect 35820 21428 35918 21664
rect 36154 21428 36252 21664
rect 36488 21428 36586 21664
rect 36822 21428 36920 21664
rect 37156 21428 37254 21664
rect 37490 21428 37588 21664
rect 37824 21428 37922 21664
rect 38158 21428 38256 21664
rect 38492 21428 38590 21664
rect 38826 21428 38924 21664
rect 39160 21428 39258 21664
rect 39494 21428 39592 21664
rect 39828 21428 40000 21664
rect 35157 21342 40000 21428
rect 35157 21106 35250 21342
rect 35486 21106 35584 21342
rect 35820 21106 35918 21342
rect 36154 21106 36252 21342
rect 36488 21106 36586 21342
rect 36822 21106 36920 21342
rect 37156 21106 37254 21342
rect 37490 21106 37588 21342
rect 37824 21106 37922 21342
rect 38158 21106 38256 21342
rect 38492 21106 38590 21342
rect 38826 21106 38924 21342
rect 39160 21106 39258 21342
rect 39494 21106 39592 21342
rect 39828 21106 40000 21342
rect 35157 21020 40000 21106
rect 35157 20784 35250 21020
rect 35486 20784 35584 21020
rect 35820 20784 35918 21020
rect 36154 20784 36252 21020
rect 36488 20784 36586 21020
rect 36822 20784 36920 21020
rect 37156 20784 37254 21020
rect 37490 20784 37588 21020
rect 37824 20784 37922 21020
rect 38158 20784 38256 21020
rect 38492 20784 38590 21020
rect 38826 20784 38924 21020
rect 39160 20784 39258 21020
rect 39494 20784 39592 21020
rect 39828 20784 40000 21020
rect 35157 20698 40000 20784
rect 35157 20462 35250 20698
rect 35486 20462 35584 20698
rect 35820 20462 35918 20698
rect 36154 20462 36252 20698
rect 36488 20462 36586 20698
rect 36822 20462 36920 20698
rect 37156 20462 37254 20698
rect 37490 20462 37588 20698
rect 37824 20462 37922 20698
rect 38158 20462 38256 20698
rect 38492 20462 38590 20698
rect 38826 20462 38924 20698
rect 39160 20462 39258 20698
rect 39494 20462 39592 20698
rect 39828 20462 40000 20698
rect 35157 20376 40000 20462
rect 35157 20140 35250 20376
rect 35486 20140 35584 20376
rect 35820 20140 35918 20376
rect 36154 20140 36252 20376
rect 36488 20140 36586 20376
rect 36822 20140 36920 20376
rect 37156 20140 37254 20376
rect 37490 20140 37588 20376
rect 37824 20140 37922 20376
rect 38158 20140 38256 20376
rect 38492 20140 38590 20376
rect 38826 20140 38924 20376
rect 39160 20140 39258 20376
rect 39494 20140 39592 20376
rect 39828 20140 40000 20376
rect 35157 20054 40000 20140
rect 35157 19818 35250 20054
rect 35486 19818 35584 20054
rect 35820 19818 35918 20054
rect 36154 19818 36252 20054
rect 36488 19818 36586 20054
rect 36822 19818 36920 20054
rect 37156 19818 37254 20054
rect 37490 19818 37588 20054
rect 37824 19818 37922 20054
rect 38158 19818 38256 20054
rect 38492 19818 38590 20054
rect 38826 19818 38924 20054
rect 39160 19818 39258 20054
rect 39494 19818 39592 20054
rect 39828 19818 40000 20054
rect 35157 19732 40000 19818
rect 0 19560 7767 19730
tri 7767 19560 7937 19730 sw
rect 0 19536 7937 19560
rect 0 19300 529 19536
rect 765 19300 863 19536
rect 1099 19300 1197 19536
rect 1433 19300 1531 19536
rect 1767 19300 1865 19536
rect 2101 19300 2199 19536
rect 2435 19300 2533 19536
rect 2769 19300 2867 19536
rect 3103 19300 3201 19536
rect 3437 19300 3535 19536
rect 3771 19300 3869 19536
rect 4105 19300 4203 19536
rect 4439 19300 4537 19536
rect 4773 19300 4871 19536
rect 5107 19300 5205 19536
rect 5441 19300 5538 19536
rect 5774 19300 5871 19536
rect 6107 19300 6204 19536
rect 6440 19300 6537 19536
rect 6773 19300 6870 19536
rect 7106 19300 7203 19536
rect 7439 19300 7536 19536
rect 7772 19300 7937 19536
rect 0 19204 7937 19300
rect 0 18968 529 19204
rect 765 18968 863 19204
rect 1099 18968 1197 19204
rect 1433 18968 1531 19204
rect 1767 18968 1865 19204
rect 2101 18968 2199 19204
rect 2435 18968 2533 19204
rect 2769 18968 2867 19204
rect 3103 18968 3201 19204
rect 3437 18968 3535 19204
rect 3771 18968 3869 19204
rect 4105 18968 4203 19204
rect 4439 18968 4537 19204
rect 4773 18968 4871 19204
rect 5107 18968 5205 19204
rect 5441 18968 5538 19204
rect 5774 18968 5871 19204
rect 6107 18968 6204 19204
rect 6440 18968 6537 19204
rect 6773 18968 6870 19204
rect 7106 18968 7203 19204
rect 7439 18968 7536 19204
rect 7772 18968 7937 19204
rect 0 18944 7937 18968
tri 7937 18944 8553 19560 sw
rect 35157 19496 35250 19732
rect 35486 19496 35584 19732
rect 35820 19496 35918 19732
rect 36154 19496 36252 19732
rect 36488 19496 36586 19732
rect 36822 19496 36920 19732
rect 37156 19496 37254 19732
rect 37490 19496 37588 19732
rect 37824 19496 37922 19732
rect 38158 19496 38256 19732
rect 38492 19496 38590 19732
rect 38826 19496 38924 19732
rect 39160 19496 39258 19732
rect 39494 19496 39592 19732
rect 39828 19496 40000 19732
rect 35157 19410 40000 19496
rect 35157 19174 35250 19410
rect 35486 19174 35584 19410
rect 35820 19174 35918 19410
rect 36154 19174 36252 19410
rect 36488 19174 36586 19410
rect 36822 19174 36920 19410
rect 37156 19174 37254 19410
rect 37490 19174 37588 19410
rect 37824 19174 37922 19410
rect 38158 19174 38256 19410
rect 38492 19174 38590 19410
rect 38826 19174 38924 19410
rect 39160 19174 39258 19410
rect 39494 19174 39592 19410
rect 39828 19174 40000 19410
rect 35157 19088 40000 19174
rect 0 18920 8553 18944
rect 0 18872 8138 18920
rect 0 18636 529 18872
rect 765 18636 863 18872
rect 1099 18636 1197 18872
rect 1433 18636 1531 18872
rect 1767 18636 1865 18872
rect 2101 18636 2199 18872
rect 2435 18636 2533 18872
rect 2769 18636 2867 18872
rect 3103 18636 3201 18872
rect 3437 18636 3535 18872
rect 3771 18636 3869 18872
rect 4105 18636 4203 18872
rect 4439 18636 4537 18872
rect 4773 18636 4871 18872
rect 5107 18636 5205 18872
rect 5441 18636 5538 18872
rect 5774 18636 5871 18872
rect 6107 18636 6204 18872
rect 6440 18636 6537 18872
rect 6773 18636 6870 18872
rect 7106 18636 7203 18872
rect 7439 18636 7536 18872
rect 7772 18684 8138 18872
rect 8374 18684 8553 18920
rect 7772 18636 8553 18684
rect 0 18596 8553 18636
rect 0 18540 8138 18596
rect 0 18304 529 18540
rect 765 18304 863 18540
rect 1099 18304 1197 18540
rect 1433 18304 1531 18540
rect 1767 18304 1865 18540
rect 2101 18304 2199 18540
rect 2435 18304 2533 18540
rect 2769 18304 2867 18540
rect 3103 18304 3201 18540
rect 3437 18304 3535 18540
rect 3771 18304 3869 18540
rect 4105 18304 4203 18540
rect 4439 18304 4537 18540
rect 4773 18304 4871 18540
rect 5107 18304 5205 18540
rect 5441 18304 5538 18540
rect 5774 18304 5871 18540
rect 6107 18304 6204 18540
rect 6440 18304 6537 18540
rect 6773 18304 6870 18540
rect 7106 18304 7203 18540
rect 7439 18304 7536 18540
rect 7772 18360 8138 18540
rect 8374 18360 8553 18596
rect 7772 18304 8553 18360
rect 0 18272 8553 18304
rect 0 18208 8138 18272
rect 0 17972 529 18208
rect 765 17972 863 18208
rect 1099 17972 1197 18208
rect 1433 17972 1531 18208
rect 1767 17972 1865 18208
rect 2101 17972 2199 18208
rect 2435 17972 2533 18208
rect 2769 17972 2867 18208
rect 3103 17972 3201 18208
rect 3437 17972 3535 18208
rect 3771 17972 3869 18208
rect 4105 17972 4203 18208
rect 4439 17972 4537 18208
rect 4773 17972 4871 18208
rect 5107 17972 5205 18208
rect 5441 17972 5538 18208
rect 5774 17972 5871 18208
rect 6107 17972 6204 18208
rect 6440 17972 6537 18208
rect 6773 17972 6870 18208
rect 7106 17972 7203 18208
rect 7439 17972 7536 18208
rect 7772 18036 8138 18208
rect 8374 18247 8553 18272
tri 8553 18247 9250 18944 sw
rect 35157 18852 35250 19088
rect 35486 18852 35584 19088
rect 35820 18852 35918 19088
rect 36154 18852 36252 19088
rect 36488 18852 36586 19088
rect 36822 18852 36920 19088
rect 37156 18852 37254 19088
rect 37490 18852 37588 19088
rect 37824 18852 37922 19088
rect 38158 18852 38256 19088
rect 38492 18852 38590 19088
rect 38826 18852 38924 19088
rect 39160 18852 39258 19088
rect 39494 18852 39592 19088
rect 39828 18852 40000 19088
rect 35157 18766 40000 18852
rect 35157 18530 35250 18766
rect 35486 18530 35584 18766
rect 35820 18530 35918 18766
rect 36154 18530 36252 18766
rect 36488 18530 36586 18766
rect 36822 18530 36920 18766
rect 37156 18530 37254 18766
rect 37490 18530 37588 18766
rect 37824 18530 37922 18766
rect 38158 18530 38256 18766
rect 38492 18530 38590 18766
rect 38826 18530 38924 18766
rect 39160 18530 39258 18766
rect 39494 18530 39592 18766
rect 39828 18530 40000 18766
rect 35157 18444 40000 18530
rect 8374 18223 9250 18247
rect 8374 18036 8835 18223
rect 7772 17987 8835 18036
rect 9071 17987 9250 18223
rect 7772 17972 9250 17987
rect 0 17948 9250 17972
rect 0 17876 8138 17948
rect 0 17640 529 17876
rect 765 17640 863 17876
rect 1099 17640 1197 17876
rect 1433 17640 1531 17876
rect 1767 17640 1865 17876
rect 2101 17640 2199 17876
rect 2435 17640 2533 17876
rect 2769 17640 2867 17876
rect 3103 17640 3201 17876
rect 3437 17640 3535 17876
rect 3771 17640 3869 17876
rect 4105 17640 4203 17876
rect 4439 17640 4537 17876
rect 4773 17640 4871 17876
rect 5107 17640 5205 17876
rect 5441 17640 5538 17876
rect 5774 17640 5871 17876
rect 6107 17640 6204 17876
rect 6440 17640 6537 17876
rect 6773 17640 6870 17876
rect 7106 17640 7203 17876
rect 7439 17640 7536 17876
rect 7772 17712 8138 17876
rect 8374 17899 9250 17948
rect 8374 17712 8835 17899
rect 7772 17663 8835 17712
rect 9071 17663 9250 17899
rect 7772 17640 9250 17663
rect 0 17624 9250 17640
rect 0 17544 8138 17624
rect 0 17308 529 17544
rect 765 17308 863 17544
rect 1099 17308 1197 17544
rect 1433 17308 1531 17544
rect 1767 17308 1865 17544
rect 2101 17308 2199 17544
rect 2435 17308 2533 17544
rect 2769 17308 2867 17544
rect 3103 17308 3201 17544
rect 3437 17308 3535 17544
rect 3771 17308 3869 17544
rect 4105 17308 4203 17544
rect 4439 17308 4537 17544
rect 4773 17308 4871 17544
rect 5107 17308 5205 17544
rect 5441 17308 5538 17544
rect 5774 17308 5871 17544
rect 6107 17308 6204 17544
rect 6440 17308 6537 17544
rect 6773 17308 6870 17544
rect 7106 17308 7203 17544
rect 7439 17308 7536 17544
rect 7772 17388 8138 17544
rect 8374 17588 9250 17624
tri 9250 17588 9909 18247 sw
rect 35157 18208 35250 18444
rect 35486 18208 35584 18444
rect 35820 18208 35918 18444
rect 36154 18208 36252 18444
rect 36488 18208 36586 18444
rect 36822 18208 36920 18444
rect 37156 18208 37254 18444
rect 37490 18208 37588 18444
rect 37824 18208 37922 18444
rect 38158 18208 38256 18444
rect 38492 18208 38590 18444
rect 38826 18208 38924 18444
rect 39160 18208 39258 18444
rect 39494 18208 39592 18444
rect 39828 18208 40000 18444
rect 35157 18122 40000 18208
rect 35157 17886 35250 18122
rect 35486 17886 35584 18122
rect 35820 17886 35918 18122
rect 36154 17886 36252 18122
rect 36488 17886 36586 18122
rect 36822 17886 36920 18122
rect 37156 17886 37254 18122
rect 37490 17886 37588 18122
rect 37824 17886 37922 18122
rect 38158 17886 38256 18122
rect 38492 17886 38590 18122
rect 38826 17886 38924 18122
rect 39160 17886 39258 18122
rect 39494 17886 39592 18122
rect 39828 17886 40000 18122
rect 35157 17800 40000 17886
rect 8374 17575 9909 17588
rect 8374 17388 8835 17575
rect 7772 17339 8835 17388
rect 9071 17564 9909 17575
rect 9071 17339 9494 17564
rect 7772 17328 9494 17339
rect 9730 17328 9909 17564
rect 7772 17308 9909 17328
rect 0 17300 9909 17308
rect 0 17212 8138 17300
rect 0 16976 529 17212
rect 765 16976 863 17212
rect 1099 16976 1197 17212
rect 1433 16976 1531 17212
rect 1767 16976 1865 17212
rect 2101 16976 2199 17212
rect 2435 16976 2533 17212
rect 2769 16976 2867 17212
rect 3103 16976 3201 17212
rect 3437 16976 3535 17212
rect 3771 16976 3869 17212
rect 4105 16976 4203 17212
rect 4439 16976 4537 17212
rect 4773 16976 4871 17212
rect 5107 16976 5205 17212
rect 5441 16976 5538 17212
rect 5774 16976 5871 17212
rect 6107 16976 6204 17212
rect 6440 16976 6537 17212
rect 6773 16976 6870 17212
rect 7106 16976 7203 17212
rect 7439 16976 7536 17212
rect 7772 17064 8138 17212
rect 8374 17251 9909 17300
rect 8374 17064 8835 17251
rect 7772 17015 8835 17064
rect 9071 17240 9909 17251
rect 9071 17015 9494 17240
rect 7772 17004 9494 17015
rect 9730 17004 9909 17240
rect 7772 16976 9909 17004
rect 0 16880 8138 16976
rect 0 16644 529 16880
rect 765 16644 863 16880
rect 1099 16644 1197 16880
rect 1433 16644 1531 16880
rect 1767 16644 1865 16880
rect 2101 16644 2199 16880
rect 2435 16644 2533 16880
rect 2769 16644 2867 16880
rect 3103 16644 3201 16880
rect 3437 16644 3535 16880
rect 3771 16644 3869 16880
rect 4105 16644 4203 16880
rect 4439 16644 4537 16880
rect 4773 16644 4871 16880
rect 5107 16644 5205 16880
rect 5441 16644 5538 16880
rect 5774 16644 5871 16880
rect 6107 16644 6204 16880
rect 6440 16644 6537 16880
rect 6773 16644 6870 16880
rect 7106 16644 7203 16880
rect 7439 16644 7536 16880
rect 7772 16740 8138 16880
rect 8374 16927 9909 16976
rect 8374 16740 8835 16927
rect 7772 16691 8835 16740
rect 9071 16916 9909 16927
rect 9071 16691 9494 16916
rect 7772 16680 9494 16691
rect 9730 16891 9909 16916
tri 9909 16891 10606 17588 sw
rect 35157 17564 35250 17800
rect 35486 17564 35584 17800
rect 35820 17564 35918 17800
rect 36154 17564 36252 17800
rect 36488 17564 36586 17800
rect 36822 17564 36920 17800
rect 37156 17564 37254 17800
rect 37490 17564 37588 17800
rect 37824 17564 37922 17800
rect 38158 17564 38256 17800
rect 38492 17564 38590 17800
rect 38826 17564 38924 17800
rect 39160 17564 39258 17800
rect 39494 17564 39592 17800
rect 39828 17564 40000 17800
rect 35157 17478 40000 17564
rect 35157 17242 35250 17478
rect 35486 17242 35584 17478
rect 35820 17242 35918 17478
rect 36154 17242 36252 17478
rect 36488 17242 36586 17478
rect 36822 17242 36920 17478
rect 37156 17242 37254 17478
rect 37490 17242 37588 17478
rect 37824 17242 37922 17478
rect 38158 17242 38256 17478
rect 38492 17242 38590 17478
rect 38826 17242 38924 17478
rect 39160 17242 39258 17478
rect 39494 17242 39592 17478
rect 39828 17242 40000 17478
rect 35157 17156 40000 17242
rect 35157 16920 35250 17156
rect 35486 16920 35584 17156
rect 35820 16920 35918 17156
rect 36154 16920 36252 17156
rect 36488 16920 36586 17156
rect 36822 16920 36920 17156
rect 37156 16920 37254 17156
rect 37490 16920 37588 17156
rect 37824 16920 37922 17156
rect 38158 16920 38256 17156
rect 38492 16920 38590 17156
rect 38826 16920 38924 17156
rect 39160 16920 39258 17156
rect 39494 16920 39592 17156
rect 39828 16920 40000 17156
rect 9730 16867 10606 16891
rect 9730 16680 10191 16867
rect 7772 16652 10191 16680
rect 7772 16644 8138 16652
rect 0 16548 8138 16644
rect 0 16312 529 16548
rect 765 16312 863 16548
rect 1099 16312 1197 16548
rect 1433 16312 1531 16548
rect 1767 16312 1865 16548
rect 2101 16312 2199 16548
rect 2435 16312 2533 16548
rect 2769 16312 2867 16548
rect 3103 16312 3201 16548
rect 3437 16312 3535 16548
rect 3771 16312 3869 16548
rect 4105 16312 4203 16548
rect 4439 16312 4537 16548
rect 4773 16312 4871 16548
rect 5107 16312 5205 16548
rect 5441 16312 5538 16548
rect 5774 16312 5871 16548
rect 6107 16312 6204 16548
rect 6440 16312 6537 16548
rect 6773 16312 6870 16548
rect 7106 16312 7203 16548
rect 7439 16312 7536 16548
rect 7772 16416 8138 16548
rect 8374 16631 10191 16652
rect 10427 16631 10606 16867
rect 8374 16603 10606 16631
rect 8374 16416 8835 16603
rect 7772 16367 8835 16416
rect 9071 16592 10606 16603
rect 9071 16367 9494 16592
rect 7772 16356 9494 16367
rect 9730 16543 10606 16592
rect 9730 16356 10191 16543
rect 7772 16328 10191 16356
rect 7772 16312 8138 16328
rect 0 16216 8138 16312
rect 0 15980 529 16216
rect 765 15980 863 16216
rect 1099 15980 1197 16216
rect 1433 15980 1531 16216
rect 1767 15980 1865 16216
rect 2101 15980 2199 16216
rect 2435 15980 2533 16216
rect 2769 15980 2867 16216
rect 3103 15980 3201 16216
rect 3437 15980 3535 16216
rect 3771 15980 3869 16216
rect 4105 15980 4203 16216
rect 4439 15980 4537 16216
rect 4773 15980 4871 16216
rect 5107 15980 5205 16216
rect 5441 15980 5538 16216
rect 5774 15980 5871 16216
rect 6107 15980 6204 16216
rect 6440 15980 6537 16216
rect 6773 15980 6870 16216
rect 7106 15980 7203 16216
rect 7439 15980 7536 16216
rect 7772 16092 8138 16216
rect 8374 16307 10191 16328
rect 10427 16307 10606 16543
rect 8374 16279 10606 16307
rect 8374 16092 8835 16279
rect 7772 16043 8835 16092
rect 9071 16268 10606 16279
rect 9071 16043 9494 16268
rect 7772 16032 9494 16043
rect 9730 16219 10606 16268
rect 9730 16032 10191 16219
rect 7772 16004 10191 16032
rect 7772 15980 8138 16004
rect 0 15884 8138 15980
rect 0 15648 529 15884
rect 765 15648 863 15884
rect 1099 15648 1197 15884
rect 1433 15648 1531 15884
rect 1767 15648 1865 15884
rect 2101 15648 2199 15884
rect 2435 15648 2533 15884
rect 2769 15648 2867 15884
rect 3103 15648 3201 15884
rect 3437 15648 3535 15884
rect 3771 15648 3869 15884
rect 4105 15648 4203 15884
rect 4439 15648 4537 15884
rect 4773 15648 4871 15884
rect 5107 15648 5205 15884
rect 5441 15648 5538 15884
rect 5774 15648 5871 15884
rect 6107 15648 6204 15884
rect 6440 15648 6537 15884
rect 6773 15648 6870 15884
rect 7106 15648 7203 15884
rect 7439 15648 7536 15884
rect 7772 15768 8138 15884
rect 8374 15983 10191 16004
rect 10427 16212 10606 16219
tri 10606 16212 11285 16891 sw
rect 35157 16834 40000 16920
rect 35157 16598 35250 16834
rect 35486 16598 35584 16834
rect 35820 16598 35918 16834
rect 36154 16598 36252 16834
rect 36488 16598 36586 16834
rect 36822 16598 36920 16834
rect 37156 16598 37254 16834
rect 37490 16598 37588 16834
rect 37824 16598 37922 16834
rect 38158 16598 38256 16834
rect 38492 16598 38590 16834
rect 38826 16598 38924 16834
rect 39160 16598 39258 16834
rect 39494 16598 39592 16834
rect 39828 16598 40000 16834
rect 35157 16512 40000 16598
rect 35157 16276 35250 16512
rect 35486 16276 35584 16512
rect 35820 16276 35918 16512
rect 36154 16276 36252 16512
rect 36488 16276 36586 16512
rect 36822 16276 36920 16512
rect 37156 16276 37254 16512
rect 37490 16276 37588 16512
rect 37824 16276 37922 16512
rect 38158 16276 38256 16512
rect 38492 16276 38590 16512
rect 38826 16276 38924 16512
rect 39160 16276 39258 16512
rect 39494 16276 39592 16512
rect 39828 16276 40000 16512
rect 10427 16188 11285 16212
rect 10427 15983 10870 16188
rect 8374 15955 10870 15983
rect 8374 15768 8835 15955
rect 7772 15719 8835 15768
rect 9071 15952 10870 15955
rect 11106 15952 11285 16188
rect 9071 15944 11285 15952
rect 9071 15719 9494 15944
rect 7772 15708 9494 15719
rect 9730 15895 11285 15944
rect 9730 15708 10191 15895
rect 7772 15680 10191 15708
rect 7772 15648 8138 15680
rect 0 15552 8138 15648
rect 0 15316 529 15552
rect 765 15316 863 15552
rect 1099 15316 1197 15552
rect 1433 15316 1531 15552
rect 1767 15316 1865 15552
rect 2101 15316 2199 15552
rect 2435 15316 2533 15552
rect 2769 15316 2867 15552
rect 3103 15316 3201 15552
rect 3437 15316 3535 15552
rect 3771 15316 3869 15552
rect 4105 15316 4203 15552
rect 4439 15316 4537 15552
rect 4773 15316 4871 15552
rect 5107 15316 5205 15552
rect 5441 15316 5538 15552
rect 5774 15316 5871 15552
rect 6107 15316 6204 15552
rect 6440 15316 6537 15552
rect 6773 15316 6870 15552
rect 7106 15316 7203 15552
rect 7439 15316 7536 15552
rect 7772 15444 8138 15552
rect 8374 15659 10191 15680
rect 10427 15864 11285 15895
rect 10427 15659 10870 15864
rect 8374 15631 10870 15659
rect 8374 15444 8835 15631
rect 7772 15395 8835 15444
rect 9071 15628 10870 15631
rect 11106 15628 11285 15864
rect 9071 15620 11285 15628
rect 9071 15395 9494 15620
rect 7772 15384 9494 15395
rect 9730 15571 11285 15620
rect 9730 15384 10191 15571
rect 7772 15356 10191 15384
rect 7772 15316 8138 15356
rect 0 15220 8138 15316
rect 0 14984 529 15220
rect 765 14984 863 15220
rect 1099 14984 1197 15220
rect 1433 14984 1531 15220
rect 1767 14984 1865 15220
rect 2101 14984 2199 15220
rect 2435 14984 2533 15220
rect 2769 14984 2867 15220
rect 3103 14984 3201 15220
rect 3437 14984 3535 15220
rect 3771 14984 3869 15220
rect 4105 14984 4203 15220
rect 4439 14984 4537 15220
rect 4773 14984 4871 15220
rect 5107 14984 5205 15220
rect 5441 14984 5538 15220
rect 5774 14984 5871 15220
rect 6107 14984 6204 15220
rect 6440 14984 6537 15220
rect 6773 14984 6870 15220
rect 7106 14984 7203 15220
rect 7439 14984 7536 15220
rect 7772 15120 8138 15220
rect 8374 15335 10191 15356
rect 10427 15540 11285 15571
rect 10427 15335 10870 15540
rect 8374 15307 10870 15335
rect 8374 15120 8835 15307
rect 7772 15071 8835 15120
rect 9071 15304 10870 15307
rect 11106 15515 11285 15540
tri 11285 15515 11982 16212 sw
rect 35157 16190 40000 16276
rect 35157 15954 35250 16190
rect 35486 15954 35584 16190
rect 35820 15954 35918 16190
rect 36154 15954 36252 16190
rect 36488 15954 36586 16190
rect 36822 15954 36920 16190
rect 37156 15954 37254 16190
rect 37490 15954 37588 16190
rect 37824 15954 37922 16190
rect 38158 15954 38256 16190
rect 38492 15954 38590 16190
rect 38826 15954 38924 16190
rect 39160 15954 39258 16190
rect 39494 15954 39592 16190
rect 39828 15954 40000 16190
rect 35157 15868 40000 15954
rect 35157 15632 35250 15868
rect 35486 15632 35584 15868
rect 35820 15632 35918 15868
rect 36154 15632 36252 15868
rect 36488 15632 36586 15868
rect 36822 15632 36920 15868
rect 37156 15632 37254 15868
rect 37490 15632 37588 15868
rect 37824 15632 37922 15868
rect 38158 15632 38256 15868
rect 38492 15632 38590 15868
rect 38826 15632 38924 15868
rect 39160 15632 39258 15868
rect 39494 15632 39592 15868
rect 39828 15632 40000 15868
rect 35157 15546 40000 15632
rect 11106 15491 11982 15515
rect 11106 15304 11567 15491
rect 9071 15296 11567 15304
rect 9071 15071 9494 15296
rect 7772 15060 9494 15071
rect 9730 15255 11567 15296
rect 11803 15255 11982 15491
rect 9730 15247 11982 15255
rect 9730 15060 10191 15247
rect 7772 15032 10191 15060
rect 7772 14984 8138 15032
rect 0 14796 8138 14984
rect 8374 15011 10191 15032
rect 10427 15216 11982 15247
rect 10427 15011 10870 15216
rect 8374 14983 10870 15011
rect 8374 14796 8835 14983
rect 0 14747 8835 14796
rect 9071 14980 10870 14983
rect 11106 15167 11982 15216
rect 11106 14980 11567 15167
rect 9071 14972 11567 14980
rect 9071 14747 9494 14972
rect 0 14740 9494 14747
tri 5739 14420 6059 14740 ne
rect 6059 14736 9494 14740
rect 9730 14931 11567 14972
rect 11803 14931 11982 15167
rect 9730 14923 11982 14931
rect 9730 14736 10191 14923
rect 6059 14708 10191 14736
rect 6059 14472 8138 14708
rect 8374 14687 10191 14708
rect 10427 14892 11982 14923
rect 10427 14687 10870 14892
rect 8374 14659 10870 14687
rect 8374 14472 8835 14659
rect 6059 14423 8835 14472
rect 9071 14656 10870 14659
rect 11106 14856 11982 14892
tri 11982 14856 12641 15515 sw
rect 35157 15310 35250 15546
rect 35486 15310 35584 15546
rect 35820 15310 35918 15546
rect 36154 15310 36252 15546
rect 36488 15310 36586 15546
rect 36822 15310 36920 15546
rect 37156 15310 37254 15546
rect 37490 15310 37588 15546
rect 37824 15310 37922 15546
rect 38158 15310 38256 15546
rect 38492 15310 38590 15546
rect 38826 15310 38924 15546
rect 39160 15310 39258 15546
rect 39494 15310 39592 15546
rect 39828 15310 40000 15546
rect 35157 15224 40000 15310
rect 35157 14988 35250 15224
rect 35486 14988 35584 15224
rect 35820 14988 35918 15224
rect 36154 14988 36252 15224
rect 36488 14988 36586 15224
rect 36822 14988 36920 15224
rect 37156 14988 37254 15224
rect 37490 14988 37588 15224
rect 37824 14988 37922 15224
rect 38158 14988 38256 15224
rect 38492 14988 38590 15224
rect 38826 14988 38924 15224
rect 39160 14988 39258 15224
rect 39494 14988 39592 15224
rect 39828 14988 40000 15224
rect 35157 14902 40000 14988
rect 11106 14843 12641 14856
rect 11106 14656 11567 14843
rect 9071 14648 11567 14656
rect 9071 14423 9494 14648
rect 6059 14420 9494 14423
rect 0 14390 5606 14420
rect 0 14154 296 14390
rect 532 14154 627 14390
rect 863 14154 958 14390
rect 1194 14154 1289 14390
rect 1525 14154 1620 14390
rect 1856 14154 1951 14390
rect 2187 14154 2282 14390
rect 2518 14154 2613 14390
rect 2849 14154 2944 14390
rect 3180 14154 3275 14390
rect 3511 14154 3606 14390
rect 3842 14154 3936 14390
rect 4172 14154 4266 14390
rect 4502 14154 4596 14390
rect 4832 14154 4926 14390
rect 5162 14154 5256 14390
rect 5492 14287 5606 14390
tri 5606 14287 5739 14420 sw
tri 6059 14287 6192 14420 ne
rect 6192 14412 9494 14420
rect 9730 14607 11567 14648
rect 11803 14832 12641 14843
rect 11803 14607 12226 14832
rect 9730 14599 12226 14607
rect 9730 14412 10191 14599
rect 6192 14384 10191 14412
rect 6192 14287 8138 14384
rect 5492 14154 5739 14287
rect 0 14116 5739 14154
tri 5739 14116 5910 14287 sw
tri 6192 14116 6363 14287 ne
rect 6363 14148 8138 14287
rect 8374 14363 10191 14384
rect 10427 14596 12226 14599
rect 12462 14740 12641 14832
tri 12641 14740 12757 14856 sw
rect 12462 14596 12757 14740
rect 10427 14568 12757 14596
rect 10427 14363 10870 14568
rect 8374 14335 10870 14363
rect 8374 14148 8835 14335
rect 6363 14116 8835 14148
rect 0 14092 5910 14116
rect 0 13856 5581 14092
rect 5817 14023 5910 14092
tri 5910 14023 6003 14116 sw
tri 6363 14023 6456 14116 ne
rect 6456 14099 8835 14116
rect 9071 14332 10870 14335
rect 11106 14519 12757 14568
rect 11106 14332 11567 14519
rect 9071 14324 11567 14332
rect 9071 14099 9494 14324
rect 6456 14088 9494 14099
rect 9730 14283 11567 14324
rect 11803 14508 12757 14519
rect 11803 14283 12226 14508
rect 9730 14275 12226 14283
rect 9730 14088 10191 14275
rect 6456 14060 10191 14088
rect 6456 14023 8138 14060
rect 5817 13856 6003 14023
rect 0 13836 6003 13856
rect 0 13600 296 13836
rect 532 13600 627 13836
rect 863 13600 958 13836
rect 1194 13600 1289 13836
rect 1525 13600 1620 13836
rect 1856 13600 1951 13836
rect 2187 13600 2282 13836
rect 2518 13600 2613 13836
rect 2849 13600 2944 13836
rect 3180 13600 3275 13836
rect 3511 13600 3606 13836
rect 3842 13600 3936 13836
rect 4172 13600 4266 13836
rect 4502 13600 4596 13836
rect 4832 13600 4926 13836
rect 5162 13600 5256 13836
rect 5492 13712 6003 13836
tri 6003 13712 6314 14023 sw
tri 6456 13712 6767 14023 ne
rect 6767 13824 8138 14023
rect 8374 14039 10191 14060
rect 10427 14272 12226 14275
rect 12462 14272 12757 14508
rect 10427 14244 12757 14272
rect 10427 14039 10870 14244
rect 8374 14011 10870 14039
rect 8374 13824 8835 14011
rect 6767 13775 8835 13824
rect 9071 14008 10870 14011
rect 11106 14195 12757 14244
rect 11106 14008 11567 14195
rect 9071 14000 11567 14008
rect 9071 13775 9494 14000
rect 6767 13764 9494 13775
rect 9730 13959 11567 14000
rect 11803 14184 12757 14195
rect 11803 13959 12226 14184
rect 9730 13951 12226 13959
rect 9730 13764 10191 13951
rect 6767 13736 10191 13764
rect 6767 13712 8138 13736
rect 5492 13688 6314 13712
rect 5492 13600 5985 13688
rect 0 13570 5985 13600
tri 5253 13285 5538 13570 ne
rect 5538 13545 5985 13570
rect 5538 13309 5581 13545
rect 5817 13452 5985 13545
rect 6221 13570 6314 13688
tri 6314 13570 6456 13712 sw
tri 6767 13570 6909 13712 ne
rect 6909 13570 8138 13712
rect 6221 13452 6456 13570
rect 5817 13309 6456 13452
rect 5538 13306 6456 13309
tri 6456 13306 6720 13570 sw
tri 6909 13306 7173 13570 ne
rect 7173 13500 8138 13570
rect 8374 13715 10191 13736
rect 10427 13948 12226 13951
rect 12462 14159 12757 14184
tri 12757 14159 13338 14740 sw
rect 35157 14666 35250 14902
rect 35486 14666 35584 14902
rect 35820 14666 35918 14902
rect 36154 14666 36252 14902
rect 36488 14666 36586 14902
rect 36822 14666 36920 14902
rect 37156 14666 37254 14902
rect 37490 14666 37588 14902
rect 37824 14666 37922 14902
rect 38158 14666 38256 14902
rect 38492 14666 38590 14902
rect 38826 14666 38924 14902
rect 39160 14666 39258 14902
rect 39494 14666 39592 14902
rect 39828 14666 40000 14902
rect 35157 14580 40000 14666
rect 35157 14344 35250 14580
rect 35486 14344 35584 14580
rect 35820 14344 35918 14580
rect 36154 14344 36252 14580
rect 36488 14344 36586 14580
rect 36822 14344 36920 14580
rect 37156 14344 37254 14580
rect 37490 14344 37588 14580
rect 37824 14344 37922 14580
rect 38158 14344 38256 14580
rect 38492 14344 38590 14580
rect 38826 14344 38924 14580
rect 39160 14344 39258 14580
rect 39494 14344 39592 14580
rect 39828 14344 40000 14580
rect 35157 14258 40000 14344
rect 12462 14135 13338 14159
rect 12462 13948 12923 14135
rect 10427 13920 12923 13948
rect 10427 13715 10870 13920
rect 8374 13687 10870 13715
rect 8374 13500 8835 13687
rect 7173 13451 8835 13500
rect 9071 13684 10870 13687
rect 11106 13899 12923 13920
rect 13159 13899 13338 14135
rect 11106 13871 13338 13899
rect 11106 13684 11567 13871
rect 9071 13676 11567 13684
rect 9071 13451 9494 13676
rect 7173 13440 9494 13451
rect 9730 13635 11567 13676
rect 11803 13860 13338 13871
rect 11803 13635 12226 13860
rect 9730 13627 12226 13635
rect 9730 13440 10191 13627
rect 7173 13412 10191 13440
rect 7173 13306 8138 13412
rect 5538 13285 6720 13306
tri 5538 13250 5573 13285 ne
rect 5573 13282 6720 13285
rect 5573 13250 6391 13282
rect 0 13239 5118 13250
tri 5118 13239 5129 13250 sw
tri 5573 13239 5584 13250 ne
rect 5584 13239 6391 13250
rect 0 13215 5129 13239
rect 0 12979 325 13215
rect 561 12979 830 13215
rect 1066 12979 1335 13215
rect 1571 12979 1840 13215
rect 2076 12979 2345 13215
rect 2581 12979 2850 13215
rect 3086 12979 3354 13215
rect 3590 12979 3858 13215
rect 4094 12979 4362 13215
rect 4598 12979 4866 13215
rect 5102 13115 5129 13215
tri 5129 13115 5253 13239 sw
tri 5584 13115 5708 13239 ne
rect 5708 13141 6391 13239
rect 5708 13115 5985 13141
rect 5102 12979 5253 13115
rect 0 12866 5253 12979
tri 5253 12866 5502 13115 sw
tri 5708 13084 5739 13115 ne
rect 5739 13084 5985 13115
tri 5739 12881 5942 13084 ne
rect 5942 12905 5985 13084
rect 6221 13046 6391 13141
rect 6627 13117 6720 13282
tri 6720 13117 6909 13306 sw
tri 7173 13117 7362 13306 ne
rect 7362 13176 8138 13306
rect 8374 13391 10191 13412
rect 10427 13624 12226 13627
rect 12462 13811 13338 13860
rect 12462 13624 12923 13811
rect 10427 13596 12923 13624
rect 10427 13391 10870 13596
rect 8374 13363 10870 13391
rect 8374 13176 8835 13363
rect 7362 13127 8835 13176
rect 9071 13360 10870 13363
rect 11106 13575 12923 13596
rect 13159 13575 13338 13811
rect 11106 13547 13338 13575
rect 11106 13360 11567 13547
rect 9071 13352 11567 13360
rect 9071 13127 9494 13352
rect 7362 13117 9494 13127
rect 6627 13046 6909 13117
rect 6221 12905 6909 13046
rect 5942 12902 6909 12905
tri 6909 12902 7124 13117 sw
tri 7362 12902 7577 13117 ne
rect 7577 13116 9494 13117
rect 9730 13311 11567 13352
rect 11803 13536 13338 13547
rect 11803 13311 12226 13536
rect 9730 13303 12226 13311
rect 9730 13116 10191 13303
rect 7577 13088 10191 13116
rect 7577 12902 8138 13088
rect 5942 12881 7124 12902
tri 5942 12866 5957 12881 ne
rect 5957 12878 7124 12881
rect 5957 12866 6795 12878
rect 0 12855 5502 12866
tri 5502 12855 5513 12866 sw
tri 5957 12855 5968 12866 ne
rect 5968 12855 6795 12866
rect 0 12842 5513 12855
rect 0 12677 5220 12842
rect 0 12441 325 12677
rect 561 12441 830 12677
rect 1066 12441 1335 12677
rect 1571 12441 1840 12677
rect 2076 12441 2345 12677
rect 2581 12441 2850 12677
rect 3086 12441 3354 12677
rect 3590 12441 3858 12677
rect 4094 12441 4362 12677
rect 4598 12441 4866 12677
rect 5102 12606 5220 12677
rect 5456 12629 5513 12842
tri 5513 12629 5739 12855 sw
tri 5968 12629 6194 12855 ne
rect 6194 12735 6795 12855
rect 6194 12629 6391 12735
rect 5456 12606 5739 12629
rect 5102 12502 5739 12606
tri 5739 12502 5866 12629 sw
tri 6194 12502 6321 12629 ne
rect 6321 12502 6391 12629
rect 5102 12478 5866 12502
rect 5102 12441 5581 12478
rect 0 12400 5581 12441
tri 4764 12367 4797 12400 ne
rect 4797 12367 5581 12400
tri 4797 12080 5084 12367 ne
rect 5084 12295 5581 12367
rect 5084 12080 5220 12295
rect 0 11627 4631 12080
tri 4631 11627 5084 12080 sw
tri 5084 12035 5129 12080 ne
rect 5129 12059 5220 12080
rect 5456 12242 5581 12295
rect 5817 12400 5866 12478
tri 5866 12400 5968 12502 sw
tri 6321 12475 6348 12502 ne
rect 6348 12499 6391 12502
rect 6627 12642 6795 12735
rect 7031 12820 7124 12878
tri 7124 12820 7206 12902 sw
tri 7577 12820 7659 12902 ne
rect 7659 12852 8138 12902
rect 8374 13067 10191 13088
rect 10427 13300 12226 13303
rect 12462 13535 13338 13536
tri 13338 13535 13962 14159 sw
rect 35157 14022 35250 14258
rect 35486 14022 35584 14258
rect 35820 14022 35918 14258
rect 36154 14022 36252 14258
rect 36488 14022 36586 14258
rect 36822 14022 36920 14258
rect 37156 14022 37254 14258
rect 37490 14022 37588 14258
rect 37824 14022 37922 14258
rect 38158 14022 38256 14258
rect 38492 14022 38590 14258
rect 38826 14022 38924 14258
rect 39160 14022 39258 14258
rect 39494 14022 39592 14258
rect 39828 14022 40000 14258
rect 35157 13936 40000 14022
rect 35157 13700 35250 13936
rect 35486 13700 35584 13936
rect 35820 13700 35918 13936
rect 36154 13700 36252 13936
rect 36488 13700 36586 13936
rect 36822 13700 36920 13936
rect 37156 13700 37254 13936
rect 37490 13700 37588 13936
rect 37824 13700 37922 13936
rect 38158 13700 38256 13936
rect 38492 13700 38590 13936
rect 38826 13700 38924 13936
rect 39160 13700 39258 13936
rect 39494 13700 39592 13936
rect 39828 13700 40000 13936
rect 35157 13614 40000 13700
rect 12462 13511 13962 13535
rect 12462 13487 13547 13511
rect 12462 13300 12923 13487
rect 10427 13272 12923 13300
rect 10427 13067 10870 13272
rect 8374 13039 10870 13067
rect 8374 12852 8835 13039
rect 7659 12820 8835 12852
rect 7031 12642 7206 12820
rect 6627 12503 7206 12642
tri 7206 12503 7523 12820 sw
tri 7659 12503 7976 12820 ne
rect 7976 12803 8835 12820
rect 9071 13036 10870 13039
rect 11106 13251 12923 13272
rect 13159 13275 13547 13487
rect 13783 13275 13962 13511
rect 13159 13251 13962 13275
rect 11106 13223 13962 13251
rect 11106 13036 11567 13223
rect 9071 13028 11567 13036
rect 9071 12803 9494 13028
rect 7976 12792 9494 12803
rect 9730 12987 11567 13028
rect 11803 13212 13962 13223
rect 11803 12987 12226 13212
rect 9730 12979 12226 12987
rect 9730 12792 10191 12979
rect 7976 12763 10191 12792
rect 7976 12527 8138 12763
rect 8374 12743 10191 12763
rect 10427 12976 12226 12979
rect 12462 13187 13962 13212
rect 12462 13163 13547 13187
rect 12462 12976 12923 13163
rect 10427 12948 12923 12976
rect 10427 12743 10870 12948
rect 8374 12715 10870 12743
rect 8374 12527 8835 12715
rect 7976 12503 8835 12527
rect 6627 12499 7523 12503
rect 6348 12479 7523 12499
rect 6348 12475 7194 12479
tri 6348 12400 6423 12475 ne
rect 6423 12400 7194 12475
rect 5817 12367 5968 12400
tri 5968 12367 6001 12400 sw
tri 6423 12367 6456 12400 ne
rect 6456 12367 7194 12400
rect 5817 12242 6001 12367
rect 5456 12098 6001 12242
tri 6001 12098 6270 12367 sw
tri 6456 12098 6725 12367 ne
rect 6725 12331 7194 12367
rect 6725 12098 6795 12331
rect 5456 12080 6270 12098
tri 6270 12080 6288 12098 sw
tri 6725 12080 6743 12098 ne
rect 6743 12095 6795 12098
rect 7031 12243 7194 12331
rect 7430 12367 7523 12479
tri 7523 12367 7659 12503 sw
tri 7976 12367 8112 12503 ne
rect 8112 12479 8835 12503
rect 9071 12712 10870 12715
rect 11106 12927 12923 12948
rect 13159 12951 13547 13163
rect 13783 12951 13962 13187
rect 13159 12927 13962 12951
rect 11106 12899 13962 12927
rect 11106 12712 11567 12899
rect 9071 12704 11567 12712
rect 9071 12479 9494 12704
rect 8112 12468 9494 12479
rect 9730 12663 11567 12704
rect 11803 12888 13962 12899
rect 11803 12663 12226 12888
rect 9730 12655 12226 12663
rect 9730 12468 10191 12655
rect 8112 12419 10191 12468
rect 10427 12652 12226 12655
rect 12462 12863 13962 12888
rect 12462 12839 13547 12863
rect 12462 12652 12923 12839
rect 10427 12624 12923 12652
rect 10427 12419 10870 12624
rect 8112 12391 10870 12419
rect 8112 12367 8835 12391
rect 7430 12243 7659 12367
rect 7031 12099 7659 12243
tri 7659 12099 7927 12367 sw
tri 8112 12099 8380 12367 ne
rect 8380 12155 8835 12367
rect 9071 12388 10870 12391
rect 11106 12603 12923 12624
rect 13159 12627 13547 12839
rect 13783 12838 13962 12863
tri 13962 12838 14659 13535 sw
rect 35157 13378 35250 13614
rect 35486 13378 35584 13614
rect 35820 13378 35918 13614
rect 36154 13378 36252 13614
rect 36488 13378 36586 13614
rect 36822 13378 36920 13614
rect 37156 13378 37254 13614
rect 37490 13378 37588 13614
rect 37824 13378 37922 13614
rect 38158 13378 38256 13614
rect 38492 13378 38590 13614
rect 38826 13378 38924 13614
rect 39160 13378 39258 13614
rect 39494 13378 39592 13614
rect 39828 13378 40000 13614
rect 35157 13292 40000 13378
rect 35157 13056 35250 13292
rect 35486 13056 35584 13292
rect 35820 13056 35918 13292
rect 36154 13056 36252 13292
rect 36488 13056 36586 13292
rect 36822 13056 36920 13292
rect 37156 13056 37254 13292
rect 37490 13056 37588 13292
rect 37824 13056 37922 13292
rect 38158 13056 38256 13292
rect 38492 13056 38590 13292
rect 38826 13056 38924 13292
rect 39160 13056 39258 13292
rect 39494 13056 39592 13292
rect 39828 13056 40000 13292
rect 35157 12970 40000 13056
rect 13783 12814 14659 12838
rect 13783 12627 14244 12814
rect 13159 12603 14244 12627
rect 11106 12578 14244 12603
rect 14480 12578 14659 12814
rect 11106 12575 14659 12578
rect 11106 12388 11567 12575
rect 9071 12380 11567 12388
rect 9071 12155 9494 12380
rect 8380 12144 9494 12155
rect 9730 12339 11567 12380
rect 11803 12564 14659 12575
rect 11803 12339 12226 12564
rect 9730 12331 12226 12339
rect 9730 12144 10191 12331
rect 8380 12099 10191 12144
rect 7031 12095 7927 12099
rect 6743 12080 7927 12095
rect 5456 12074 6288 12080
rect 5456 12059 5985 12074
rect 5129 12035 5985 12059
tri 5129 11627 5537 12035 ne
rect 5537 11931 5985 12035
rect 5537 11695 5581 11931
rect 5817 11838 5985 11931
rect 6221 11937 6288 12074
tri 6288 11937 6431 12080 sw
tri 6743 12071 6752 12080 ne
rect 6752 12075 7927 12080
rect 6752 12071 7598 12075
tri 6752 11937 6886 12071 ne
rect 6886 11937 7598 12071
rect 6221 11912 6431 11937
tri 6431 11912 6456 11937 sw
tri 6886 11912 6911 11937 ne
rect 6911 11932 7598 11937
rect 6911 11912 7194 11932
rect 6221 11838 6456 11912
rect 5817 11695 6456 11838
rect 5537 11692 6456 11695
tri 6456 11692 6676 11912 sw
tri 6911 11692 7131 11912 ne
rect 7131 11696 7194 11912
rect 7430 11839 7598 11932
rect 7834 11914 7927 12075
tri 7927 11914 8112 12099 sw
tri 8380 11914 8565 12099 ne
rect 8565 12095 10191 12099
rect 10427 12328 12226 12331
rect 12462 12539 14659 12564
rect 12462 12515 13547 12539
rect 12462 12328 12923 12515
rect 10427 12300 12923 12328
rect 10427 12095 10870 12300
rect 8565 12066 10870 12095
rect 8565 11914 8835 12066
rect 7834 11839 8112 11914
rect 7430 11696 8112 11839
rect 7131 11692 8112 11696
rect 5537 11668 6676 11692
rect 5537 11627 6391 11668
rect 0 11425 5084 11627
tri 5084 11425 5286 11627 sw
tri 5537 11425 5739 11627 ne
rect 5739 11527 6391 11627
rect 5739 11425 5985 11527
rect 0 11196 5286 11425
tri 5286 11196 5515 11425 sw
tri 5739 11267 5897 11425 ne
rect 5897 11291 5985 11425
rect 6221 11432 6391 11527
rect 6627 11651 6676 11668
tri 6676 11651 6717 11692 sw
tri 7131 11672 7151 11692 ne
rect 7151 11688 8112 11692
tri 8112 11688 8338 11914 sw
tri 8565 11806 8673 11914 ne
rect 8673 11830 8835 11914
rect 9071 12064 10870 12066
rect 11106 12279 12923 12300
rect 13159 12303 13547 12515
rect 13783 12492 14659 12539
rect 13783 12303 14244 12492
rect 13159 12279 14244 12303
rect 11106 12256 14244 12279
rect 14480 12256 14659 12492
rect 11106 12251 14659 12256
rect 11106 12064 11567 12251
rect 9071 12056 11567 12064
rect 9071 11830 9494 12056
rect 8673 11820 9494 11830
rect 9730 12015 11567 12056
rect 11803 12240 14659 12251
rect 11803 12015 12226 12240
rect 9730 12007 12226 12015
rect 9730 11820 10191 12007
rect 8673 11806 10191 11820
tri 8673 11688 8791 11806 ne
rect 8791 11771 10191 11806
rect 10427 12004 12226 12007
rect 12462 12215 14659 12240
rect 12462 12191 13547 12215
rect 12462 12004 12923 12191
rect 10427 11976 12923 12004
rect 10427 11771 10870 11976
rect 8791 11740 10870 11771
rect 11106 11955 12923 11976
rect 13159 11979 13547 12191
rect 13783 12179 14659 12215
tri 14659 12179 15318 12838 sw
rect 35157 12734 35250 12970
rect 35486 12734 35584 12970
rect 35820 12734 35918 12970
rect 36154 12734 36252 12970
rect 36488 12734 36586 12970
rect 36822 12734 36920 12970
rect 37156 12734 37254 12970
rect 37490 12734 37588 12970
rect 37824 12734 37922 12970
rect 38158 12734 38256 12970
rect 38492 12734 38590 12970
rect 38826 12734 38924 12970
rect 39160 12734 39258 12970
rect 39494 12734 39592 12970
rect 39828 12734 40000 12970
rect 35157 12648 40000 12734
rect 35157 12412 35250 12648
rect 35486 12412 35584 12648
rect 35820 12412 35918 12648
rect 36154 12412 36252 12648
rect 36488 12412 36586 12648
rect 36822 12412 36920 12648
rect 37156 12412 37254 12648
rect 37490 12412 37588 12648
rect 37824 12412 37922 12648
rect 38158 12412 38256 12648
rect 38492 12412 38590 12648
rect 38826 12412 38924 12648
rect 39160 12412 39258 12648
rect 39494 12412 39592 12648
rect 39828 12412 40000 12648
rect 35157 12326 40000 12412
rect 13783 12170 15318 12179
rect 13783 11979 14244 12170
rect 13159 11955 14244 11979
rect 11106 11934 14244 11955
rect 14480 12155 15318 12170
rect 14480 11934 14903 12155
rect 11106 11927 14903 11934
rect 11106 11740 11567 11927
rect 8791 11732 11567 11740
rect 8791 11688 9494 11732
rect 7151 11672 8338 11688
tri 7151 11651 7172 11672 ne
rect 7172 11664 8338 11672
rect 7172 11651 8009 11664
rect 6627 11432 6717 11651
rect 6221 11291 6717 11432
rect 5897 11286 6717 11291
tri 6717 11286 7082 11651 sw
tri 7172 11286 7537 11651 ne
rect 7537 11528 8009 11651
rect 7537 11292 7598 11528
rect 7834 11428 8009 11528
rect 8245 11617 8338 11664
tri 8338 11617 8409 11688 sw
tri 8791 11617 8862 11688 ne
rect 8862 11617 9494 11688
rect 8245 11428 8409 11617
rect 7834 11292 8409 11428
rect 7537 11286 8409 11292
rect 5897 11267 7082 11286
tri 5897 11196 5968 11267 ne
rect 5968 11262 7082 11267
rect 5968 11196 6800 11262
rect 0 11164 5515 11196
tri 5515 11164 5547 11196 sw
tri 5968 11164 6000 11196 ne
rect 6000 11164 6800 11196
rect 0 10733 5547 11164
tri 5547 10733 5978 11164 sw
tri 6000 10861 6303 11164 ne
rect 6303 11121 6800 11164
rect 6303 10885 6391 11121
rect 6627 11026 6800 11121
rect 7036 11196 7082 11262
tri 7082 11196 7172 11286 sw
tri 7537 11268 7555 11286 ne
rect 7555 11284 8409 11286
tri 8409 11284 8742 11617 sw
tri 8862 11284 9195 11617 ne
rect 9195 11496 9494 11617
rect 9730 11691 11567 11732
rect 11803 11919 14903 11927
rect 15139 11919 15318 12155
rect 11803 11916 15318 11919
rect 11803 11691 12226 11916
rect 9730 11683 12226 11691
rect 9730 11496 10191 11683
rect 9195 11447 10191 11496
rect 10427 11680 12226 11683
rect 12462 11891 15318 11916
rect 12462 11867 13547 11891
rect 12462 11680 12923 11867
rect 10427 11652 12923 11680
rect 10427 11447 10870 11652
rect 9195 11416 10870 11447
rect 11106 11631 12923 11652
rect 13159 11655 13547 11867
rect 13783 11848 15318 11891
rect 13783 11655 14244 11848
rect 13159 11631 14244 11655
rect 11106 11612 14244 11631
rect 14480 11834 15318 11848
rect 14480 11612 14903 11834
rect 11106 11603 14903 11612
rect 11106 11416 11567 11603
rect 9195 11407 11567 11416
rect 9195 11284 9494 11407
rect 7555 11268 8742 11284
tri 7555 11196 7627 11268 ne
rect 7627 11260 8742 11268
rect 7627 11196 8413 11260
rect 7036 11164 7172 11196
tri 7172 11164 7204 11196 sw
tri 7627 11164 7659 11196 ne
rect 7659 11164 8413 11196
rect 7036 11026 7204 11164
rect 6627 10922 7204 11026
tri 7204 10922 7446 11164 sw
tri 7659 10922 7901 11164 ne
rect 7901 11117 8413 11164
rect 7901 10922 8009 11117
rect 6627 10898 7446 10922
rect 6627 10885 7161 10898
rect 6303 10861 7161 10885
tri 6303 10733 6431 10861 ne
rect 6431 10733 7161 10861
rect 0 10280 5978 10733
tri 5978 10280 6431 10733 sw
tri 6431 10455 6709 10733 ne
rect 6709 10715 7161 10733
rect 6709 10479 6800 10715
rect 7036 10662 7161 10715
rect 7397 10709 7446 10898
tri 7446 10709 7659 10922 sw
tri 7901 10857 7966 10922 ne
rect 7966 10881 8009 10922
rect 8245 11024 8413 11117
rect 8649 11164 8742 11260
tri 8742 11164 8862 11284 sw
tri 9195 11164 9315 11284 ne
rect 9315 11171 9494 11284
rect 9730 11367 11567 11407
rect 11803 11598 14903 11603
rect 15139 11598 15318 11834
rect 11803 11592 15318 11598
rect 11803 11367 12226 11592
rect 9730 11359 12226 11367
rect 9730 11171 10191 11359
rect 9315 11164 10191 11171
rect 8649 11024 8862 11164
rect 8245 10885 8862 11024
tri 8862 10885 9141 11164 sw
tri 9315 11147 9332 11164 ne
rect 9332 11147 10191 11164
tri 9332 10885 9594 11147 ne
rect 9594 11123 10191 11147
rect 10427 11356 12226 11359
rect 12462 11567 15318 11592
rect 12462 11543 13547 11567
rect 12462 11356 12923 11543
rect 10427 11328 12923 11356
rect 10427 11123 10870 11328
rect 9594 11092 10870 11123
rect 11106 11307 12923 11328
rect 13159 11331 13547 11543
rect 13783 11526 15318 11567
rect 13783 11331 14244 11526
rect 13159 11307 14244 11331
rect 11106 11290 14244 11307
rect 14480 11513 15318 11526
rect 14480 11290 14903 11513
rect 11106 11279 14903 11290
rect 11106 11092 11567 11279
rect 9594 11043 11567 11092
rect 11803 11277 14903 11279
rect 15139 11482 15318 11513
tri 15318 11482 16015 12179 sw
rect 35157 12090 35250 12326
rect 35486 12090 35584 12326
rect 35820 12090 35918 12326
rect 36154 12090 36252 12326
rect 36488 12090 36586 12326
rect 36822 12090 36920 12326
rect 37156 12090 37254 12326
rect 37490 12090 37588 12326
rect 37824 12090 37922 12326
rect 38158 12090 38256 12326
rect 38492 12090 38590 12326
rect 38826 12090 38924 12326
rect 39160 12090 39258 12326
rect 39494 12090 39592 12326
rect 39828 12090 40000 12326
rect 35157 12004 40000 12090
rect 35157 11768 35250 12004
rect 35486 11768 35584 12004
rect 35820 11768 35918 12004
rect 36154 11768 36252 12004
rect 36488 11768 36586 12004
rect 36822 11768 36920 12004
rect 37156 11768 37254 12004
rect 37490 11768 37588 12004
rect 37824 11768 37922 12004
rect 38158 11768 38256 12004
rect 38492 11768 38590 12004
rect 38826 11768 38924 12004
rect 39160 11768 39258 12004
rect 39494 11768 39592 12004
rect 39828 11768 40000 12004
rect 35157 11682 40000 11768
rect 15139 11458 16015 11482
rect 15139 11277 15600 11458
rect 11803 11268 15600 11277
rect 11803 11043 12226 11268
rect 9594 11035 12226 11043
rect 9594 10885 10191 11035
rect 8245 10881 9141 10885
rect 7966 10861 9141 10881
rect 7966 10857 8812 10861
tri 7966 10709 8114 10857 ne
rect 8114 10713 8812 10857
rect 8114 10709 8413 10713
rect 7397 10662 7659 10709
rect 7036 10518 7659 10662
tri 7659 10518 7850 10709 sw
tri 8114 10518 8305 10709 ne
rect 8305 10518 8413 10709
rect 7036 10494 7850 10518
rect 7036 10479 7565 10494
rect 6709 10455 7565 10479
tri 6709 10280 6884 10455 ne
rect 6884 10351 7565 10455
rect 6884 10280 7161 10351
tri 3887 9992 4175 10280 ne
rect 4175 9992 6431 10280
tri 6431 9992 6719 10280 sw
tri 6884 10091 7073 10280 ne
rect 7073 10115 7161 10280
rect 7397 10258 7565 10351
rect 7801 10447 7850 10494
tri 7850 10447 7921 10518 sw
tri 8305 10447 8376 10518 ne
rect 8376 10477 8413 10518
rect 8649 10625 8812 10713
rect 9048 10711 9141 10861
tri 9141 10711 9315 10885 sw
tri 9594 10711 9768 10885 ne
rect 9768 10799 10191 10885
rect 10427 11032 12226 11035
rect 12462 11243 15600 11268
rect 12462 11219 13547 11243
rect 12462 11032 12923 11219
rect 10427 11004 12923 11032
rect 10427 10799 10870 11004
rect 9768 10768 10870 10799
rect 11106 10983 12923 11004
rect 13159 11007 13547 11219
rect 13783 11222 15600 11243
rect 15836 11222 16015 11458
rect 13783 11204 16015 11222
rect 13783 11007 14244 11204
rect 13159 10983 14244 11007
rect 11106 10968 14244 10983
rect 14480 11192 16015 11204
rect 14480 10968 14903 11192
rect 11106 10956 14903 10968
rect 15139 11127 16015 11192
rect 15139 10956 15600 11127
rect 11106 10955 15600 10956
rect 11106 10768 11567 10955
rect 9768 10719 11567 10768
rect 11803 10944 15600 10955
rect 11803 10719 12226 10944
rect 9768 10711 12226 10719
rect 9048 10625 9315 10711
rect 8649 10481 9315 10625
tri 9315 10481 9545 10711 sw
tri 9768 10481 9998 10711 ne
rect 9998 10710 12226 10711
rect 9998 10481 10191 10710
rect 8649 10477 9545 10481
rect 8376 10457 9545 10477
rect 8376 10447 9216 10457
rect 7801 10280 7921 10447
tri 7921 10280 8088 10447 sw
tri 8376 10280 8543 10447 ne
rect 8543 10314 9216 10447
rect 8543 10280 8812 10314
rect 7801 10258 8088 10280
rect 7397 10115 8088 10258
rect 7073 10112 8088 10115
tri 8088 10112 8256 10280 sw
tri 8543 10112 8711 10280 ne
rect 8711 10112 8812 10280
rect 7073 10091 8256 10112
tri 7073 9992 7172 10091 ne
rect 7172 10088 8256 10091
rect 7172 9992 7971 10088
tri 4175 9960 4207 9992 ne
rect 4207 9960 6719 9992
tri 6719 9960 6751 9992 sw
tri 7172 9960 7204 9992 ne
rect 7204 9960 7971 9992
rect 0 9944 3754 9960
tri 3754 9944 3770 9960 sw
tri 4207 9944 4223 9960 ne
rect 4223 9944 6751 9960
rect 0 9920 3770 9944
rect 0 9684 295 9920
rect 531 9684 830 9920
rect 1066 9684 1365 9920
rect 1601 9684 1900 9920
rect 2136 9684 2434 9920
rect 2670 9684 2968 9920
rect 3204 9684 3502 9920
rect 3738 9827 3770 9920
tri 3770 9827 3887 9944 sw
tri 4223 9827 4340 9944 ne
rect 4340 9827 6751 9944
rect 3738 9684 3887 9827
rect 0 9565 3887 9684
tri 3887 9565 4149 9827 sw
tri 4340 9565 4602 9827 ne
rect 4602 9565 6751 9827
rect 0 9541 4149 9565
rect 0 9346 3820 9541
rect 0 9110 295 9346
rect 531 9110 830 9346
rect 1066 9110 1365 9346
rect 1601 9110 1900 9346
rect 2136 9110 2434 9346
rect 2670 9110 2968 9346
rect 3204 9110 3502 9346
rect 3738 9305 3820 9346
rect 4056 9523 4149 9541
tri 4149 9523 4191 9565 sw
tri 4602 9523 4644 9565 ne
rect 4644 9523 6751 9565
rect 4056 9305 4191 9523
rect 3738 9206 4191 9305
tri 4191 9206 4508 9523 sw
tri 4644 9206 4961 9523 ne
rect 4961 9507 6751 9523
tri 6751 9507 7204 9960 sw
tri 7204 9687 7477 9960 ne
rect 7477 9947 7971 9960
rect 7477 9711 7565 9947
rect 7801 9852 7971 9947
rect 8207 9992 8256 10088
tri 8256 9992 8376 10112 sw
tri 8711 10054 8769 10112 ne
rect 8769 10078 8812 10112
rect 9048 10221 9216 10314
rect 9452 10414 9545 10457
tri 9545 10414 9612 10481 sw
tri 9998 10414 10065 10481 ne
rect 10065 10474 10191 10481
rect 10427 10708 12226 10710
rect 12462 10919 15600 10944
rect 12462 10895 13547 10919
rect 12462 10708 12923 10895
rect 10427 10680 12923 10708
rect 10427 10474 10870 10680
rect 10065 10444 10870 10474
rect 11106 10659 12923 10680
rect 13159 10683 13547 10895
rect 13783 10891 15600 10919
rect 15836 11121 16015 11127
tri 16015 11121 16376 11482 sw
rect 35157 11446 35250 11682
rect 35486 11446 35584 11682
rect 35820 11446 35918 11682
rect 36154 11446 36252 11682
rect 36488 11446 36586 11682
rect 36822 11446 36920 11682
rect 37156 11446 37254 11682
rect 37490 11446 37588 11682
rect 37824 11446 37922 11682
rect 38158 11446 38256 11682
rect 38492 11446 38590 11682
rect 38826 11446 38924 11682
rect 39160 11446 39258 11682
rect 39494 11446 39592 11682
rect 39828 11446 40000 11682
rect 35157 11360 40000 11446
rect 35157 11124 35250 11360
rect 35486 11124 35584 11360
rect 35820 11124 35918 11360
rect 36154 11124 36252 11360
rect 36488 11124 36586 11360
rect 36822 11124 36920 11360
rect 37156 11124 37254 11360
rect 37490 11124 37588 11360
rect 37824 11124 37922 11360
rect 38158 11124 38256 11360
rect 38492 11124 38590 11360
rect 38826 11124 38924 11360
rect 39160 11124 39258 11360
rect 39494 11124 39592 11360
rect 39828 11124 40000 11360
rect 15836 11097 16386 11121
rect 15836 10891 16073 11097
rect 13783 10882 16073 10891
rect 13783 10683 14244 10882
rect 13159 10659 14244 10683
rect 11106 10646 14244 10659
rect 14480 10871 16073 10882
rect 14480 10646 14903 10871
rect 11106 10635 14903 10646
rect 15139 10861 16073 10871
rect 16309 10861 16386 11097
rect 15139 10796 16386 10861
rect 15139 10635 15600 10796
rect 11106 10631 15600 10635
rect 11106 10444 11567 10631
rect 10065 10414 11567 10444
rect 9452 10221 9612 10414
rect 9048 10078 9612 10221
rect 8769 10054 9612 10078
tri 8769 9992 8831 10054 ne
rect 8831 10048 9612 10054
tri 9612 10048 9978 10414 sw
tri 10065 10048 10431 10414 ne
rect 10431 10395 11567 10414
rect 11803 10620 15600 10631
rect 11803 10395 12226 10620
rect 10431 10384 12226 10395
rect 12462 10595 15600 10620
rect 12462 10571 13547 10595
rect 12462 10384 12923 10571
rect 10431 10356 12923 10384
rect 10431 10120 10870 10356
rect 11106 10335 12923 10356
rect 13159 10359 13547 10571
rect 13783 10560 15600 10595
rect 15836 10560 16386 10796
rect 13783 10359 14244 10560
rect 13159 10335 14244 10359
rect 11106 10324 14244 10335
rect 14480 10550 16386 10560
rect 14480 10324 14903 10550
rect 11106 10314 14903 10324
rect 15139 10465 16386 10550
rect 15139 10314 15600 10465
rect 11106 10307 15600 10314
rect 11106 10120 11567 10307
rect 10431 10071 11567 10120
rect 11803 10296 15600 10307
rect 11803 10071 12226 10296
rect 10431 10060 12226 10071
rect 12462 10271 15600 10296
rect 12462 10247 13547 10271
rect 12462 10060 12923 10247
rect 10431 10048 12923 10060
rect 8831 10024 9978 10048
rect 8831 9992 9649 10024
rect 8207 9961 8376 9992
tri 8376 9961 8407 9992 sw
tri 8831 9961 8862 9992 ne
rect 8862 9961 9649 9992
rect 8207 9852 8407 9961
rect 7801 9721 8407 9852
tri 8407 9721 8647 9961 sw
tri 8862 9848 8975 9961 ne
rect 8975 9910 9649 9961
rect 8975 9848 9216 9910
tri 8975 9721 9102 9848 ne
rect 9102 9721 9216 9848
rect 7801 9711 8647 9721
rect 7477 9697 8647 9711
rect 7477 9687 8365 9697
tri 7477 9507 7657 9687 ne
rect 7657 9541 8365 9687
rect 7657 9507 7971 9541
rect 4961 9206 7204 9507
rect 3738 9182 4508 9206
rect 3738 9110 4195 9182
rect 0 9070 4195 9110
tri 3390 8750 3710 9070 ne
rect 3710 8994 4195 9070
rect 3710 8758 3820 8994
rect 4056 8946 4195 8994
rect 4431 9070 4508 9182
tri 4508 9070 4644 9206 sw
tri 4961 9070 5097 9206 ne
rect 5097 9070 7204 9206
tri 7204 9070 7641 9507 sw
tri 7657 9281 7883 9507 ne
rect 7883 9305 7971 9507
rect 8207 9461 8365 9541
rect 8601 9506 8647 9697
tri 8647 9506 8862 9721 sw
tri 9102 9650 9173 9721 ne
rect 9173 9674 9216 9721
rect 9452 9788 9649 9910
rect 9885 9961 9978 10024
tri 9978 9961 10065 10048 sw
tri 10431 9961 10518 10048 ne
rect 10518 10031 12923 10048
rect 10518 9961 10870 10031
rect 9885 9788 10065 9961
rect 9452 9674 10065 9788
rect 9173 9650 10065 9674
tri 9173 9506 9317 9650 ne
rect 9317 9644 10065 9650
tri 10065 9644 10382 9961 sw
tri 10518 9771 10708 9961 ne
rect 10708 9795 10870 9961
rect 11106 10011 12923 10031
rect 13159 10035 13547 10247
rect 13783 10238 15600 10271
rect 13783 10035 14244 10238
rect 13159 10011 14244 10035
rect 11106 10002 14244 10011
rect 14480 10229 15600 10238
rect 15836 10462 16386 10465
rect 15836 10229 16073 10462
rect 14480 10002 14903 10229
rect 11106 9993 14903 10002
rect 15139 10226 16073 10229
rect 16309 10226 16386 10462
rect 15139 10202 16386 10226
tri 16386 10202 17295 11111 sw
rect 35157 11038 40000 11124
rect 35157 10802 35250 11038
rect 35486 10802 35584 11038
rect 35820 10802 35918 11038
rect 36154 10802 36252 11038
rect 36488 10802 36586 11038
rect 36822 10802 36920 11038
rect 37156 10802 37254 11038
rect 37490 10802 37588 11038
rect 37824 10802 37922 11038
rect 38158 10802 38256 11038
rect 38492 10802 38590 11038
rect 38826 10802 38924 11038
rect 39160 10802 39258 11038
rect 39494 10802 39592 11038
rect 39828 10802 40000 11038
rect 35157 10716 40000 10802
rect 35157 10480 35250 10716
rect 35486 10480 35584 10716
rect 35820 10480 35918 10716
rect 36154 10480 36252 10716
rect 36488 10480 36586 10716
rect 36822 10480 36920 10716
rect 37156 10480 37254 10716
rect 37490 10480 37588 10716
rect 37824 10480 37922 10716
rect 38158 10480 38256 10716
rect 38492 10480 38590 10716
rect 38826 10480 38924 10716
rect 39160 10480 39258 10716
rect 39494 10480 39592 10716
rect 39828 10480 40000 10716
rect 35157 10394 40000 10480
rect 15139 10192 17295 10202
tri 17295 10192 17305 10202 sw
rect 15139 10134 17305 10192
rect 15139 9993 15600 10134
rect 11106 9983 15600 9993
rect 11106 9795 11567 9983
rect 10708 9771 11567 9795
tri 10708 9644 10835 9771 ne
rect 10835 9747 11567 9771
rect 11803 9972 15600 9983
rect 11803 9747 12226 9972
rect 10835 9736 12226 9747
rect 12462 9947 15600 9972
rect 12462 9923 13547 9947
rect 12462 9736 12923 9923
rect 10835 9687 12923 9736
rect 13159 9711 13547 9923
rect 13783 9915 15600 9947
rect 13783 9711 14244 9915
rect 13159 9687 14244 9711
rect 10835 9679 14244 9687
rect 14480 9908 15600 9915
rect 14480 9679 14903 9908
rect 10835 9672 14903 9679
rect 15139 9898 15600 9908
rect 15836 10079 17305 10134
rect 15836 9898 16050 10079
rect 15139 9843 16050 9898
rect 16286 9843 16545 10079
rect 16781 9843 17039 10079
rect 17275 9843 17305 10079
rect 15139 9803 17305 9843
rect 15139 9672 15600 9803
rect 10835 9659 15600 9672
rect 10835 9644 11567 9659
rect 9317 9620 10382 9644
rect 9317 9506 10053 9620
rect 8601 9461 8862 9506
rect 8207 9393 8862 9461
tri 8862 9393 8975 9506 sw
tri 9317 9393 9430 9506 ne
rect 9430 9477 10053 9506
rect 9430 9393 9649 9477
rect 8207 9357 8975 9393
tri 8975 9357 9011 9393 sw
tri 9430 9357 9466 9393 ne
rect 9466 9357 9649 9393
rect 8207 9333 9011 9357
rect 8207 9305 8726 9333
rect 7883 9281 8726 9305
tri 7883 9070 8094 9281 ne
rect 8094 9150 8726 9281
rect 8094 9070 8365 9150
rect 4431 8946 4644 9070
rect 4056 8842 4644 8946
tri 4644 8842 4872 9070 sw
tri 5097 8842 5325 9070 ne
rect 5325 8842 7641 9070
rect 4056 8818 4872 8842
rect 4056 8758 4556 8818
rect 3710 8750 4556 8758
rect 0 8726 3257 8750
tri 3257 8726 3281 8750 sw
tri 3710 8734 3726 8750 ne
rect 3726 8734 4556 8750
tri 3726 8726 3734 8734 ne
rect 3734 8726 4556 8734
rect 0 8702 3281 8726
rect 0 8466 267 8702
rect 503 8466 816 8702
rect 1052 8466 1365 8702
rect 1601 8466 1914 8702
rect 2150 8466 2463 8702
rect 2699 8466 3012 8702
rect 3248 8617 3281 8702
tri 3281 8617 3390 8726 sw
tri 3734 8617 3843 8726 ne
rect 3843 8635 4556 8726
rect 3843 8617 4195 8635
rect 3248 8590 3390 8617
tri 3390 8590 3417 8617 sw
tri 3843 8590 3870 8617 ne
rect 3870 8590 4195 8617
rect 3248 8466 3417 8590
rect 0 8362 3417 8466
rect 0 8126 267 8362
rect 503 8126 816 8362
rect 1052 8126 1365 8362
rect 1601 8126 1914 8362
rect 2150 8126 2463 8362
rect 2699 8126 3012 8362
rect 3248 8269 3417 8362
tri 3417 8269 3738 8590 sw
tri 3870 8573 3887 8590 ne
rect 3887 8573 4195 8590
tri 3887 8375 4085 8573 ne
rect 4085 8399 4195 8573
rect 4431 8582 4556 8635
rect 4792 8617 4872 8818
tri 4872 8617 5097 8842 sw
tri 5325 8617 5550 8842 ne
rect 5550 8788 7641 8842
tri 7641 8788 7923 9070 sw
tri 8094 8890 8274 9070 ne
rect 8274 8914 8365 9070
rect 8601 9097 8726 9150
rect 8962 9243 9011 9333
tri 9011 9243 9125 9357 sw
tri 9466 9243 9580 9357 ne
rect 9580 9243 9649 9357
rect 8962 9097 9125 9243
rect 8601 8953 9125 9097
tri 9125 8953 9415 9243 sw
tri 9580 9217 9606 9243 ne
rect 9606 9241 9649 9243
rect 9885 9384 10053 9477
rect 10289 9508 10382 9620
tri 10382 9508 10518 9644 sw
tri 10835 9508 10971 9644 ne
rect 10971 9508 11567 9644
rect 10289 9384 10518 9508
rect 9885 9245 10518 9384
tri 10518 9245 10781 9508 sw
tri 10971 9245 11234 9508 ne
rect 11234 9423 11567 9508
rect 11803 9648 15600 9659
rect 11803 9423 12226 9648
rect 11234 9412 12226 9423
rect 12462 9623 15600 9648
rect 12462 9599 13547 9623
rect 12462 9412 12923 9599
rect 11234 9363 12923 9412
rect 13159 9387 13547 9599
rect 13783 9592 15600 9623
rect 13783 9387 14244 9592
rect 13159 9363 14244 9387
rect 11234 9356 14244 9363
rect 14480 9587 15600 9592
rect 14480 9356 14903 9587
rect 11234 9351 14903 9356
rect 15139 9567 15600 9587
rect 15836 9624 17305 9803
tri 17305 9624 17873 10192 sw
rect 35157 10158 35250 10394
rect 35486 10158 35584 10394
rect 35820 10158 35918 10394
rect 36154 10158 36252 10394
rect 36488 10158 36586 10394
rect 36822 10158 36920 10394
rect 37156 10158 37254 10394
rect 37490 10158 37588 10394
rect 37824 10158 37922 10394
rect 38158 10158 38256 10394
rect 38492 10158 38590 10394
rect 38826 10158 38924 10394
rect 39160 10158 39258 10394
rect 39494 10158 39592 10394
rect 39828 10158 40000 10394
rect 35157 10072 40000 10158
rect 35157 9836 35250 10072
rect 35486 9836 35584 10072
rect 35820 9836 35918 10072
rect 36154 9836 36252 10072
rect 36488 9836 36586 10072
rect 36822 9836 36920 10072
rect 37156 9836 37254 10072
rect 37490 9836 37588 10072
rect 37824 9836 37922 10072
rect 38158 9836 38256 10072
rect 38492 9836 38590 10072
rect 38826 9836 38924 10072
rect 39160 9836 39258 10072
rect 39494 9836 39592 10072
rect 39828 9836 40000 10072
rect 35157 9750 40000 9836
rect 15836 9599 17873 9624
rect 15836 9567 16065 9599
rect 15139 9471 16065 9567
rect 15139 9351 15600 9471
rect 11234 9334 15600 9351
rect 11234 9245 11567 9334
rect 9885 9241 10781 9245
rect 9606 9221 10781 9241
rect 9606 9217 10452 9221
tri 9606 8953 9870 9217 ne
rect 9870 9073 10452 9217
rect 9870 8953 10053 9073
rect 8601 8929 9415 8953
rect 8601 8914 9130 8929
rect 8274 8890 9130 8914
tri 8274 8788 8376 8890 ne
rect 8376 8788 9130 8890
rect 5550 8758 7923 8788
tri 7923 8758 7953 8788 sw
tri 8376 8758 8406 8788 ne
rect 8406 8786 9130 8788
rect 8406 8758 8726 8786
rect 5550 8617 7953 8758
rect 4792 8582 5097 8617
rect 4431 8456 5097 8582
tri 5097 8456 5258 8617 sw
tri 5550 8456 5711 8617 ne
rect 5711 8456 7953 8617
rect 4431 8432 5258 8456
rect 4431 8399 4945 8432
rect 4085 8375 4945 8399
tri 4085 8269 4191 8375 ne
rect 4191 8271 4945 8375
rect 4191 8269 4556 8271
rect 3248 8126 3738 8269
rect 0 8120 3738 8126
tri 3738 8120 3887 8269 sw
tri 4191 8120 4340 8269 ne
rect 4340 8120 4556 8269
rect 0 8100 3887 8120
tri 2987 7780 3307 8100 ne
rect 3307 7816 3887 8100
tri 3887 7816 4191 8120 sw
tri 4340 8011 4449 8120 ne
rect 4449 8035 4556 8120
rect 4792 8196 4945 8271
rect 5181 8428 5258 8432
tri 5258 8428 5286 8456 sw
tri 5711 8428 5739 8456 ne
rect 5739 8428 7953 8456
rect 5181 8196 5286 8428
rect 4792 8092 5286 8196
tri 5286 8092 5622 8428 sw
tri 5739 8092 6075 8428 ne
rect 6075 8305 7953 8428
tri 7953 8305 8406 8758 sw
tri 8406 8526 8638 8758 ne
rect 8638 8550 8726 8758
rect 8962 8693 9130 8786
rect 9366 8788 9415 8929
tri 9415 8788 9580 8953 sw
tri 9870 8813 10010 8953 ne
rect 10010 8837 10053 8953
rect 10289 8985 10452 9073
rect 10688 9211 10781 9221
tri 10781 9211 10815 9245 sw
tri 11234 9211 11268 9245 ne
rect 11268 9211 11567 9245
rect 10688 8985 10815 9211
rect 10289 8841 10815 8985
tri 10815 8841 11185 9211 sw
tri 11268 9074 11405 9211 ne
rect 11405 9098 11567 9211
rect 11803 9324 15600 9334
rect 11803 9098 12226 9324
rect 11405 9088 12226 9098
rect 12462 9299 15600 9324
rect 12462 9275 13547 9299
rect 12462 9088 12923 9275
rect 11405 9074 12923 9088
tri 11405 8841 11638 9074 ne
rect 11638 9039 12923 9074
rect 13159 9063 13547 9275
rect 13783 9269 15600 9299
rect 13783 9063 14244 9269
rect 13159 9039 14244 9063
rect 11638 9033 14244 9039
rect 14480 9266 15600 9269
rect 14480 9033 14903 9266
rect 11638 9030 14903 9033
rect 15139 9235 15600 9266
rect 15836 9363 16065 9471
rect 16301 9363 16575 9599
rect 16811 9363 17084 9599
rect 17320 9363 17593 9599
rect 17829 9363 17873 9599
rect 15836 9261 17873 9363
rect 15836 9235 16065 9261
rect 15139 9139 16065 9235
rect 15139 9030 15600 9139
rect 11638 9000 15600 9030
rect 11638 8841 12226 9000
rect 10289 8837 11185 8841
rect 10010 8817 11185 8837
rect 10010 8813 10856 8817
tri 10010 8788 10035 8813 ne
rect 10035 8788 10856 8813
rect 9366 8758 9580 8788
tri 9580 8758 9610 8788 sw
tri 10035 8758 10065 8788 ne
rect 10065 8758 10856 8788
rect 9366 8693 9610 8758
rect 8962 8550 9610 8693
rect 8638 8547 9610 8550
tri 9610 8547 9821 8758 sw
tri 10065 8547 10276 8758 ne
rect 10276 8674 10856 8758
rect 10276 8547 10452 8674
rect 8638 8526 9821 8547
tri 8638 8305 8859 8526 ne
rect 8859 8523 9821 8526
rect 8859 8382 9536 8523
rect 8859 8305 9130 8382
rect 6075 8189 8406 8305
tri 8406 8189 8522 8305 sw
tri 8859 8189 8975 8305 ne
rect 8975 8189 9130 8305
rect 6075 8092 8522 8189
rect 4792 8068 5622 8092
rect 4792 8035 5306 8068
rect 4449 8011 5306 8035
tri 4449 7816 4644 8011 ne
rect 4644 7885 5306 8011
rect 4644 7816 4945 7885
rect 3307 7780 4191 7816
tri 4191 7780 4227 7816 sw
tri 4644 7780 4680 7816 ne
rect 4680 7780 4945 7816
rect 0 7762 2854 7780
tri 2854 7762 2872 7780 sw
tri 3307 7762 3325 7780 ne
rect 3325 7762 4227 7780
rect 0 7738 2872 7762
rect 0 7502 277 7738
rect 513 7502 860 7738
rect 1096 7502 1442 7738
rect 1678 7502 2024 7738
rect 2260 7502 2606 7738
rect 2842 7670 2872 7738
tri 2872 7670 2964 7762 sw
tri 3325 7670 3417 7762 ne
rect 3417 7736 4227 7762
tri 4227 7736 4271 7780 sw
tri 4680 7736 4724 7780 ne
rect 4724 7736 4945 7780
rect 3417 7670 4271 7736
tri 4271 7670 4337 7736 sw
tri 4724 7670 4790 7736 ne
rect 4790 7670 4945 7736
rect 2842 7502 2964 7670
rect 0 7400 2964 7502
rect 0 7164 277 7400
rect 513 7164 860 7400
rect 1096 7164 1442 7400
rect 1678 7164 2024 7400
rect 2260 7164 2606 7400
rect 2842 7217 2964 7400
tri 2964 7217 3417 7670 sw
tri 3417 7217 3870 7670 ne
rect 3870 7363 4337 7670
tri 4337 7363 4644 7670 sw
tri 4790 7625 4835 7670 ne
rect 4835 7649 4945 7670
rect 5181 7832 5306 7885
rect 5542 7975 5622 8068
tri 5622 7975 5739 8092 sw
tri 6075 7975 6192 8092 ne
rect 6192 7975 8522 8092
rect 5542 7832 5739 7975
rect 5181 7816 5739 7832
tri 5739 7816 5898 7975 sw
tri 6192 7816 6351 7975 ne
rect 6351 7816 8522 7975
tri 8522 7816 8895 8189 sw
tri 8975 8122 9042 8189 ne
rect 9042 8146 9130 8189
rect 9366 8287 9536 8382
rect 9772 8303 9821 8523
tri 9821 8303 10065 8547 sw
tri 10276 8414 10409 8547 ne
rect 10409 8438 10452 8547
rect 10688 8581 10856 8674
rect 11092 8758 11185 8817
tri 11185 8758 11268 8841 sw
tri 11638 8758 11721 8841 ne
rect 11721 8764 12226 8841
rect 12462 8975 15600 9000
rect 12462 8951 13547 8975
rect 12462 8764 12923 8951
rect 11721 8758 12923 8764
rect 11092 8581 11268 8758
rect 10688 8438 11268 8581
rect 10409 8414 11268 8438
tri 10409 8303 10520 8414 ne
rect 10520 8394 11268 8414
tri 11268 8394 11632 8758 sw
tri 11721 8415 12064 8758 ne
rect 12064 8715 12923 8758
rect 13159 8739 13547 8951
rect 13783 8946 15600 8975
rect 13783 8739 14244 8946
rect 13159 8715 14244 8739
rect 12064 8710 14244 8715
rect 14480 8945 15600 8946
rect 14480 8710 14903 8945
rect 12064 8709 14903 8710
rect 15139 8903 15600 8945
rect 15836 9025 16065 9139
rect 16301 9025 16575 9261
rect 16811 9025 17084 9261
rect 17320 9025 17593 9261
rect 17829 9025 17873 9261
rect 15836 8923 17873 9025
rect 15836 8903 16065 8923
rect 15139 8807 16065 8903
rect 15139 8709 15600 8807
rect 12064 8675 15600 8709
rect 12064 8439 12226 8675
rect 12462 8651 15600 8675
rect 12462 8627 13547 8651
rect 12462 8439 12923 8627
rect 12064 8415 12923 8439
tri 12064 8394 12085 8415 ne
rect 12085 8394 12923 8415
rect 10520 8370 11632 8394
rect 10520 8303 11303 8370
rect 9772 8287 10065 8303
rect 9366 8146 10065 8287
rect 9042 8131 10065 8146
tri 10065 8131 10237 8303 sw
tri 10520 8131 10692 8303 ne
rect 10692 8270 11303 8303
rect 10692 8131 10856 8270
rect 9042 8122 10237 8131
tri 9042 7816 9348 8122 ne
rect 9348 8107 10237 8122
rect 9348 7976 9955 8107
rect 9348 7816 9536 7976
rect 5181 7736 5898 7816
tri 5898 7736 5978 7816 sw
tri 6351 7736 6431 7816 ne
rect 6431 7736 8895 7816
tri 8895 7736 8975 7816 sw
tri 9348 7736 9428 7816 ne
rect 9428 7740 9536 7816
rect 9772 7871 9955 7976
rect 10191 8039 10237 8107
tri 10237 8039 10329 8131 sw
tri 10692 8039 10784 8131 ne
rect 10784 8039 10856 8131
rect 10191 7871 10329 8039
rect 9772 7767 10329 7871
tri 10329 7767 10601 8039 sw
tri 10784 8010 10813 8039 ne
rect 10813 8034 10856 8039
rect 11092 8134 11303 8270
rect 11539 8305 11632 8370
tri 11632 8305 11721 8394 sw
tri 12085 8305 12174 8394 ne
rect 12174 8391 12923 8394
rect 13159 8415 13547 8627
rect 13783 8624 15600 8651
rect 13783 8623 14903 8624
rect 13783 8415 14244 8623
rect 13159 8391 14244 8415
rect 12174 8387 14244 8391
rect 14480 8388 14903 8623
rect 15139 8571 15600 8624
rect 15836 8687 16065 8807
rect 16301 8687 16575 8923
rect 16811 8687 17084 8923
rect 17320 8687 17593 8923
rect 17829 8687 17873 8923
rect 15836 8571 17873 8687
rect 15139 8525 17873 8571
tri 17873 8525 18972 9624 sw
rect 35157 9514 35250 9750
rect 35486 9514 35584 9750
rect 35820 9514 35918 9750
rect 36154 9514 36252 9750
rect 36488 9514 36586 9750
rect 36822 9514 36920 9750
rect 37156 9514 37254 9750
rect 37490 9514 37588 9750
rect 37824 9514 37922 9750
rect 38158 9514 38256 9750
rect 38492 9514 38590 9750
rect 38826 9514 38924 9750
rect 39160 9514 39258 9750
rect 39494 9514 39592 9750
rect 39828 9514 40000 9750
rect 35157 9428 40000 9514
rect 35157 9192 35250 9428
rect 35486 9192 35584 9428
rect 35820 9192 35918 9428
rect 36154 9192 36252 9428
rect 36488 9192 36586 9428
rect 36822 9192 36920 9428
rect 37156 9192 37254 9428
rect 37490 9192 37588 9428
rect 37824 9192 37922 9428
rect 38158 9192 38256 9428
rect 38492 9192 38590 9428
rect 38826 9192 38924 9428
rect 39160 9192 39258 9428
rect 39494 9192 39592 9428
rect 39828 9192 40000 9428
rect 35157 9106 40000 9192
rect 35157 8870 35250 9106
rect 35486 8870 35584 9106
rect 35820 8870 35918 9106
rect 36154 8870 36252 9106
rect 36488 8870 36586 9106
rect 36822 8870 36920 9106
rect 37156 8870 37254 9106
rect 37490 8870 37588 9106
rect 37824 8870 37922 9106
rect 38158 8870 38256 9106
rect 38492 8870 38590 9106
rect 38826 8870 38924 9106
rect 39160 8870 39258 9106
rect 39494 8870 39592 9106
rect 39828 8870 40000 9106
rect 35157 8784 40000 8870
rect 35157 8548 35250 8784
rect 35486 8548 35584 8784
rect 35820 8548 35918 8784
rect 36154 8548 36252 8784
rect 36488 8548 36586 8784
rect 36822 8548 36920 8784
rect 37156 8548 37254 8784
rect 37490 8548 37588 8784
rect 37824 8548 37922 8784
rect 38158 8548 38256 8784
rect 38492 8548 38590 8784
rect 38826 8548 38924 8784
rect 39160 8548 39258 8784
rect 39494 8548 39592 8784
rect 39828 8548 40000 8784
rect 15139 8501 18972 8525
rect 15139 8475 16047 8501
rect 15139 8388 15600 8475
rect 14480 8387 15600 8388
rect 12174 8327 15600 8387
rect 12174 8305 13547 8327
rect 11539 8175 11721 8305
tri 11721 8175 11851 8305 sw
tri 12174 8175 12304 8305 ne
rect 12304 8303 13547 8305
rect 12304 8175 12923 8303
rect 11539 8134 11851 8175
rect 11092 8034 11851 8134
rect 10813 8010 11851 8034
tri 10813 7767 11056 8010 ne
rect 11056 7990 11851 8010
tri 11851 7990 12036 8175 sw
tri 12304 7990 12489 8175 ne
rect 12489 8067 12923 8175
rect 13159 8091 13547 8303
rect 13783 8302 15600 8327
rect 13783 8300 14903 8302
rect 13783 8091 14244 8300
rect 13159 8067 14244 8091
rect 12489 8064 14244 8067
rect 14480 8066 14903 8300
rect 15139 8239 15600 8302
rect 15836 8265 16047 8475
rect 16283 8265 16549 8501
rect 16785 8265 17050 8501
rect 17286 8265 17551 8501
rect 17787 8265 18052 8501
rect 18288 8265 18553 8501
rect 18789 8500 18972 8501
tri 18972 8500 18997 8525 sw
rect 18789 8265 18997 8500
rect 15836 8239 18997 8265
rect 15139 8143 18997 8239
rect 15139 8066 15600 8143
rect 14480 8064 15600 8066
rect 12489 8003 15600 8064
rect 12489 7990 13547 8003
rect 11056 7966 12036 7990
rect 11056 7823 11707 7966
rect 11056 7767 11303 7823
rect 9772 7743 10601 7767
rect 9772 7740 10316 7743
rect 9428 7736 10316 7740
rect 5181 7722 5978 7736
tri 5978 7722 5992 7736 sw
tri 6431 7722 6445 7736 ne
rect 6445 7722 8975 7736
tri 8975 7722 8989 7736 sw
tri 9428 7722 9442 7736 ne
rect 9442 7722 10316 7736
rect 5181 7669 5992 7722
rect 5181 7649 5692 7669
rect 4835 7625 5692 7649
tri 4835 7363 5097 7625 ne
rect 5097 7521 5692 7625
rect 5097 7363 5306 7521
rect 3870 7217 4644 7363
rect 2842 7164 3417 7217
rect 0 7130 3417 7164
tri 3417 7130 3504 7217 sw
tri 3870 7130 3957 7217 ne
rect 3957 7130 4644 7217
tri 4644 7130 4877 7363 sw
tri 5097 7261 5199 7363 ne
rect 5199 7285 5306 7363
rect 5542 7433 5692 7521
rect 5928 7433 5992 7669
rect 5542 7334 5992 7433
tri 5992 7334 6380 7722 sw
tri 6445 7584 6583 7722 ne
rect 6583 7584 8989 7722
tri 8989 7584 9127 7722 sw
tri 9442 7716 9448 7722 ne
rect 9448 7716 10316 7722
tri 9448 7584 9580 7716 ne
rect 9580 7584 10316 7716
tri 6583 7555 6612 7584 ne
rect 6612 7555 9127 7584
tri 9127 7555 9156 7584 sw
tri 9580 7555 9609 7584 ne
rect 9609 7560 10316 7584
rect 9609 7555 9955 7560
tri 6612 7334 6833 7555 ne
rect 6833 7334 9156 7555
rect 5542 7310 6380 7334
rect 5542 7285 6067 7310
rect 5199 7261 6067 7285
tri 5199 7130 5330 7261 ne
rect 5330 7130 6067 7261
tri 2587 6810 2907 7130 ne
rect 2907 6810 3504 7130
rect 0 6749 2454 6810
rect 0 6513 320 6749
rect 556 6513 786 6749
rect 1022 6513 1252 6749
rect 1488 6513 1718 6749
rect 1954 6513 2183 6749
rect 2419 6677 2454 6749
tri 2454 6677 2587 6810 sw
tri 2907 6677 3040 6810 ne
rect 3040 6750 3504 6810
tri 3504 6750 3884 7130 sw
tri 3957 6750 4337 7130 ne
rect 4337 6750 4877 7130
tri 4877 6750 5257 7130 sw
tri 5330 6862 5598 7130 ne
rect 5598 7122 6067 7130
rect 5598 6886 5692 7122
rect 5928 7074 6067 7122
rect 6303 7283 6380 7310
tri 6380 7283 6431 7334 sw
tri 6833 7283 6884 7334 ne
rect 6884 7283 9156 7334
rect 6303 7074 6431 7283
rect 5928 7015 6431 7074
tri 6431 7015 6699 7283 sw
tri 6884 7015 7152 7283 ne
rect 7152 7102 9156 7283
tri 9156 7102 9609 7555 sw
tri 9609 7300 9864 7555 ne
rect 9864 7324 9955 7555
rect 10191 7507 10316 7560
rect 10552 7736 10601 7743
tri 10601 7736 10632 7767 sw
tri 11056 7736 11087 7767 ne
rect 11087 7736 11303 7767
rect 10552 7722 10632 7736
tri 10632 7722 10646 7736 sw
tri 11087 7722 11101 7736 ne
rect 11101 7722 11303 7736
rect 10552 7584 10646 7722
tri 10646 7584 10784 7722 sw
tri 11101 7584 11239 7722 ne
rect 11239 7587 11303 7722
rect 11539 7730 11707 7823
rect 11943 7730 12036 7966
rect 11539 7722 12036 7730
tri 12036 7722 12304 7990 sw
tri 12489 7722 12757 7990 ne
rect 12757 7978 13547 7990
rect 12757 7742 12923 7978
rect 13159 7767 13547 7978
rect 13783 7980 15600 8003
rect 13783 7977 14903 7980
rect 13783 7767 14244 7977
rect 13159 7742 14244 7767
rect 12757 7741 14244 7742
rect 14480 7744 14903 7977
rect 15139 7907 15600 7980
rect 15836 8089 18997 8143
rect 15836 7907 16047 8089
rect 15139 7853 16047 7907
rect 16283 7853 16549 8089
rect 16785 7853 17050 8089
rect 17286 7853 17551 8089
rect 17787 7853 18052 8089
rect 18288 7853 18553 8089
rect 18789 7853 18997 8089
rect 15139 7811 18997 7853
rect 15139 7744 15600 7811
rect 14480 7741 15600 7744
rect 12757 7722 15600 7741
rect 11539 7591 12304 7722
tri 12304 7591 12435 7722 sw
tri 12757 7718 12761 7722 ne
rect 12761 7718 15600 7722
tri 12761 7591 12888 7718 ne
rect 12888 7679 15600 7718
rect 12888 7591 13547 7679
rect 11539 7587 12435 7591
rect 11239 7584 12435 7587
rect 10552 7555 10784 7584
tri 10784 7555 10813 7584 sw
tri 11239 7555 11268 7584 ne
rect 11268 7567 12435 7584
rect 11268 7555 12106 7567
rect 10552 7507 10813 7555
rect 10191 7363 10813 7507
tri 10813 7363 11005 7555 sw
tri 11268 7476 11347 7555 ne
rect 11347 7476 12106 7555
tri 11347 7363 11460 7476 ne
rect 11460 7419 12106 7476
rect 11460 7363 11707 7419
rect 10191 7339 11005 7363
rect 10191 7324 10720 7339
rect 9864 7300 10720 7324
tri 9864 7102 10062 7300 ne
rect 10062 7196 10720 7300
rect 10062 7102 10316 7196
rect 7152 7015 9609 7102
tri 9609 7015 9696 7102 sw
tri 10062 7015 10149 7102 ne
rect 10149 7015 10316 7102
rect 5928 6946 6699 7015
rect 5928 6886 6428 6946
rect 5598 6862 6428 6886
tri 5598 6750 5710 6862 ne
rect 5710 6763 6428 6862
rect 5710 6750 6067 6763
rect 3040 6677 3884 6750
rect 2419 6666 2587 6677
tri 2587 6666 2598 6677 sw
tri 3040 6666 3051 6677 ne
rect 3051 6666 3884 6677
rect 2419 6513 2598 6666
rect 0 6495 2598 6513
tri 2598 6495 2769 6666 sw
tri 3051 6495 3222 6666 ne
rect 3222 6495 3884 6666
rect 0 6471 2769 6495
rect 0 6235 2506 6471
rect 2742 6235 2769 6471
rect 0 6215 2769 6235
rect 0 5979 320 6215
rect 556 5979 786 6215
rect 1022 5979 1252 6215
rect 1488 5979 1718 6215
rect 1954 5979 2183 6215
rect 2419 6213 2769 6215
tri 2769 6213 3051 6495 sw
tri 3222 6213 3504 6495 ne
rect 3504 6297 3884 6495
tri 3884 6297 4337 6750 sw
tri 4337 6562 4525 6750 ne
rect 4525 6562 5257 6750
tri 5257 6562 5445 6750 sw
tri 5710 6562 5898 6750 ne
rect 5898 6562 6067 6750
tri 4525 6297 4790 6562 ne
rect 4790 6297 5445 6562
rect 3504 6213 4337 6297
tri 4337 6213 4421 6297 sw
tri 4790 6213 4874 6297 ne
rect 4874 6213 5445 6297
tri 5445 6213 5794 6562 sw
tri 5898 6503 5957 6562 ne
rect 5957 6527 6067 6562
rect 6303 6710 6428 6763
rect 6664 6710 6699 6946
rect 6303 6584 6699 6710
tri 6699 6584 7130 7015 sw
tri 7152 6584 7583 7015 ne
rect 7583 6584 9696 7015
rect 6303 6562 7130 6584
tri 7130 6562 7152 6584 sw
tri 7583 6562 7605 6584 ne
rect 7605 6562 9696 6584
tri 9696 6562 10149 7015 sw
tri 10149 6936 10228 7015 ne
rect 10228 6960 10316 7015
rect 10552 7103 10720 7196
rect 10956 7103 11005 7339
rect 10552 7100 11005 7103
tri 11005 7100 11268 7363 sw
tri 11460 7159 11664 7363 ne
rect 11664 7183 11707 7363
rect 11943 7331 12106 7419
rect 12342 7555 12435 7567
tri 12435 7555 12471 7591 sw
tri 12888 7555 12924 7591 ne
rect 12924 7555 13547 7591
rect 12342 7331 12471 7555
rect 11943 7269 12471 7331
tri 12471 7269 12757 7555 sw
tri 12924 7269 13210 7555 ne
rect 13210 7443 13547 7555
rect 13783 7658 15600 7679
rect 13783 7654 14903 7658
rect 13783 7443 14244 7654
rect 13210 7418 14244 7443
rect 14480 7422 14903 7654
rect 15139 7575 15600 7658
rect 15836 7677 18997 7811
rect 15836 7575 16047 7677
rect 15139 7479 16047 7575
rect 15139 7422 15600 7479
rect 14480 7418 15600 7422
rect 13210 7354 15600 7418
rect 13210 7269 13547 7354
rect 11943 7189 12757 7269
tri 12757 7189 12837 7269 sw
tri 13210 7189 13290 7269 ne
rect 13290 7189 13547 7269
rect 11943 7183 12837 7189
rect 11664 7163 12837 7183
rect 11664 7159 12510 7163
tri 11664 7100 11723 7159 ne
rect 11723 7100 12510 7159
rect 10552 7021 11268 7100
tri 11268 7021 11347 7100 sw
tri 11723 7021 11802 7100 ne
rect 11802 7021 12510 7100
rect 10552 6960 11347 7021
rect 10228 6957 11347 6960
tri 11347 6957 11411 7021 sw
tri 11802 6957 11866 7021 ne
rect 11866 7020 12510 7021
rect 11866 6957 12106 7020
rect 10228 6936 11411 6957
tri 10228 6562 10602 6936 ne
rect 10602 6933 11411 6936
rect 10602 6792 11126 6933
rect 10602 6562 10720 6792
rect 6303 6560 7152 6562
rect 6303 6527 6817 6560
rect 5957 6503 6817 6527
tri 5957 6213 6247 6503 ne
rect 6247 6399 6817 6503
rect 6247 6213 6428 6399
rect 2419 6144 3051 6213
rect 2419 5979 2506 6144
rect 0 5920 2506 5979
tri 2085 5705 2300 5920 ne
rect 2300 5908 2506 5920
rect 2742 6113 3051 6144
tri 3051 6113 3151 6213 sw
tri 3504 6113 3604 6213 ne
rect 3604 6113 4421 6213
rect 2742 6089 3151 6113
rect 2742 5908 2888 6089
rect 2300 5853 2888 5908
rect 3124 5853 3151 6089
rect 2300 5816 3151 5853
rect 2300 5705 2506 5816
tri 2300 5600 2405 5705 ne
rect 2405 5600 2506 5705
rect 0 5566 1952 5600
tri 1952 5566 1986 5600 sw
tri 2405 5566 2439 5600 ne
rect 2439 5580 2506 5600
rect 2742 5762 3151 5816
rect 2742 5580 2888 5762
rect 2439 5566 2888 5580
rect 0 5551 1986 5566
tri 1986 5551 2001 5566 sw
tri 2439 5551 2454 5566 ne
rect 2454 5551 2888 5566
rect 0 5542 2001 5551
rect 0 5306 305 5542
rect 541 5306 772 5542
rect 1008 5306 1239 5542
rect 1475 5306 1706 5542
rect 1942 5306 2001 5542
rect 0 5145 2001 5306
tri 2001 5145 2407 5551 sw
tri 2454 5174 2831 5551 ne
rect 2831 5526 2888 5551
rect 3124 5760 3151 5762
tri 3151 5760 3504 6113 sw
tri 3604 5760 3957 6113 ne
rect 3957 5830 4421 6113
tri 4421 5830 4804 6213 sw
tri 4874 5830 5257 6213 ne
rect 5257 6109 5794 6213
tri 5794 6109 5898 6213 sw
tri 6247 6109 6351 6213 ne
rect 6351 6163 6428 6213
rect 6664 6324 6817 6399
rect 7053 6324 7152 6560
rect 6664 6220 7152 6324
tri 7152 6220 7494 6562 sw
tri 7605 6220 7947 6562 ne
rect 7947 6380 10149 6562
tri 10149 6380 10331 6562 sw
tri 10602 6532 10632 6562 ne
rect 10632 6556 10720 6562
rect 10956 6697 11126 6792
rect 11362 6701 11411 6933
tri 11411 6701 11667 6957 sw
tri 11866 6760 12063 6957 ne
rect 12063 6784 12106 6957
rect 12342 6927 12510 7020
rect 12746 6927 12837 7163
rect 12342 6925 12837 6927
tri 12837 6925 13101 7189 sw
tri 13290 7094 13385 7189 ne
rect 13385 7118 13547 7189
rect 13783 7336 15600 7354
rect 13783 7331 14903 7336
rect 13783 7118 14244 7331
rect 13385 7095 14244 7118
rect 14480 7100 14903 7331
rect 15139 7243 15600 7336
rect 15836 7441 16047 7479
rect 16283 7441 16549 7677
rect 16785 7441 17050 7677
rect 17286 7441 17551 7677
rect 17787 7441 18052 7677
rect 18288 7441 18553 7677
rect 18789 7441 18997 7677
rect 15836 7265 18997 7441
rect 15836 7243 16047 7265
rect 15139 7147 16047 7243
rect 15139 7100 15600 7147
rect 14480 7095 15600 7100
rect 13385 7094 15600 7095
tri 13385 6925 13554 7094 ne
rect 13554 6925 15600 7094
rect 12342 6784 13101 6925
rect 12063 6760 13101 6784
tri 12063 6701 12122 6760 ne
rect 12122 6701 13101 6760
rect 11362 6697 11667 6701
rect 10956 6556 11667 6697
rect 10632 6532 11667 6556
tri 10632 6380 10784 6532 ne
rect 10784 6386 11667 6532
rect 10784 6380 11126 6386
rect 7947 6352 10331 6380
tri 10331 6352 10359 6380 sw
tri 10784 6352 10812 6380 ne
rect 10812 6352 11126 6380
rect 7947 6220 10359 6352
rect 6664 6196 7494 6220
rect 6664 6163 7178 6196
rect 6351 6109 7178 6163
rect 5257 5830 5898 6109
tri 5898 5830 6177 6109 sw
tri 6351 6029 6431 6109 ne
rect 6431 6029 7178 6109
tri 6431 5830 6630 6029 ne
rect 6630 6013 7178 6029
rect 6630 5830 6817 6013
rect 3957 5760 4804 5830
rect 3124 5705 3504 5760
tri 3504 5705 3559 5760 sw
tri 3957 5705 4012 5760 ne
rect 4012 5705 4804 5760
rect 3124 5700 3559 5705
tri 3559 5700 3564 5705 sw
tri 4012 5700 4017 5705 ne
rect 4017 5700 4804 5705
rect 3124 5676 3564 5700
rect 3124 5526 3301 5676
rect 2831 5440 3301 5526
rect 3537 5600 3564 5676
tri 3564 5600 3664 5700 sw
tri 4017 5600 4117 5700 ne
rect 4117 5600 4804 5700
rect 3537 5440 3664 5600
rect 2831 5434 3664 5440
rect 2831 5198 2888 5434
rect 3124 5349 3664 5434
rect 3124 5198 3301 5349
rect 2831 5174 3301 5198
tri 2831 5145 2860 5174 ne
rect 2860 5145 3301 5174
rect 0 5121 2407 5145
rect 0 4980 2139 5121
rect 0 4744 305 4980
rect 541 4744 772 4980
rect 1008 4744 1239 4980
rect 1475 4744 1706 4980
rect 1942 4885 2139 4980
rect 2375 5098 2407 5121
tri 2407 5098 2454 5145 sw
tri 2860 5098 2907 5145 ne
rect 2907 5113 3301 5145
rect 3537 5318 3664 5349
tri 3664 5318 3946 5600 sw
tri 4117 5318 4399 5600 ne
rect 4399 5377 4804 5600
tri 4804 5377 5257 5830 sw
tri 5257 5377 5710 5830 ne
rect 5710 5761 6177 5830
tri 6177 5761 6246 5830 sw
tri 6630 5761 6699 5830 ne
rect 6699 5777 6817 5830
rect 7053 5960 7178 6013
rect 7414 6109 7494 6196
tri 7494 6109 7605 6220 sw
tri 7947 6109 8058 6220 ne
rect 8058 6109 10359 6220
rect 7414 5960 7605 6109
rect 7053 5830 7605 5960
tri 7605 5830 7884 6109 sw
tri 8058 5830 8337 6109 ne
rect 8337 5899 10359 6109
tri 10359 5899 10812 6352 sw
tri 10812 6126 11038 6352 ne
rect 11038 6150 11126 6352
rect 11362 6380 11667 6386
tri 11667 6380 11988 6701 sw
tri 12122 6380 12443 6701 ne
rect 12443 6616 13101 6701
rect 12443 6380 12510 6616
rect 12746 6472 13101 6616
tri 13101 6472 13554 6925 sw
tri 13554 6472 14007 6925 ne
rect 14007 6911 15600 6925
rect 15836 7029 16047 7147
rect 16283 7029 16549 7265
rect 16785 7029 17050 7265
rect 17286 7029 17551 7265
rect 17787 7029 18052 7265
rect 18288 7029 18553 7265
rect 18789 7029 18997 7265
rect 15836 6911 18997 7029
rect 14007 6853 18997 6911
rect 14007 6617 16047 6853
rect 16283 6617 16549 6853
rect 16785 6617 17050 6853
rect 17286 6617 17551 6853
rect 17787 6617 18052 6853
rect 18288 6617 18553 6853
rect 18789 6617 18997 6853
rect 14007 6489 18997 6617
rect 12746 6380 13554 6472
rect 11362 6352 11988 6380
tri 11988 6352 12016 6380 sw
tri 12443 6352 12471 6380 ne
rect 12471 6352 13554 6380
tri 13554 6352 13674 6472 sw
rect 11362 6150 12016 6352
rect 11038 6126 12016 6150
tri 11038 5899 11265 6126 ne
rect 11265 5986 12016 6126
tri 12016 5986 12382 6352 sw
tri 12471 5986 12837 6352 ne
rect 12837 6339 13674 6352
tri 13674 6339 13687 6352 sw
rect 12837 6279 13687 6339
rect 12837 6043 12869 6279
rect 13105 6043 13421 6279
rect 13657 6043 13687 6279
rect 11265 5899 12382 5986
rect 8337 5830 10812 5899
rect 7053 5788 7884 5830
rect 7053 5777 7589 5788
rect 6699 5761 7589 5777
rect 5710 5576 6246 5761
tri 6246 5576 6431 5761 sw
tri 6699 5753 6707 5761 ne
rect 6707 5753 7589 5761
tri 6707 5576 6884 5753 ne
rect 6884 5649 7589 5753
rect 6884 5576 7178 5649
rect 5710 5377 6431 5576
rect 4399 5318 5257 5377
rect 3537 5296 3946 5318
tri 3946 5296 3968 5318 sw
tri 4399 5296 4421 5318 ne
rect 4421 5296 5257 5318
tri 5257 5296 5338 5377 sw
tri 5710 5296 5791 5377 ne
rect 5791 5308 6431 5377
tri 6431 5308 6699 5576 sw
tri 6884 5308 7152 5576 ne
rect 7152 5413 7178 5576
rect 7414 5552 7589 5649
rect 7825 5552 7884 5788
rect 7414 5448 7884 5552
tri 7884 5448 8266 5830 sw
tri 8337 5497 8670 5830 ne
rect 8670 5817 10812 5830
tri 10812 5817 10894 5899 sw
tri 11265 5817 11347 5899 ne
rect 11347 5851 12382 5899
tri 12382 5851 12517 5986 sw
rect 11347 5817 12517 5851
rect 8670 5497 10894 5817
tri 10894 5497 11214 5817 sw
tri 11347 5497 11667 5817 ne
rect 11667 5812 12517 5817
rect 11667 5576 11703 5812
rect 11939 5576 12237 5812
rect 12473 5576 12517 5812
tri 8670 5448 8719 5497 ne
rect 8719 5448 11214 5497
rect 7414 5424 8266 5448
rect 7414 5413 7950 5424
rect 7152 5308 7950 5413
rect 5791 5296 6699 5308
tri 6699 5296 6711 5308 sw
tri 7152 5296 7164 5308 ne
rect 7164 5296 7950 5308
rect 3537 5294 3968 5296
rect 3537 5113 3683 5294
rect 2907 5098 3683 5113
rect 2375 4885 2454 5098
rect 1942 4794 2454 4885
rect 1942 4744 2139 4794
rect 0 4710 2139 4744
tri 1583 4390 1903 4710 ne
rect 1903 4558 2139 4710
rect 2375 4763 2454 4794
tri 2454 4763 2789 5098 sw
tri 2907 4763 3242 5098 ne
rect 3242 5058 3683 5098
rect 3919 5058 3968 5294
rect 3242 5021 3968 5058
rect 3242 4785 3301 5021
rect 3537 4967 3968 5021
rect 3537 4785 3683 4967
rect 3242 4763 3683 4785
rect 2375 4739 2789 4763
rect 2375 4558 2521 4739
rect 1903 4503 2521 4558
rect 2757 4710 2789 4739
tri 2789 4710 2842 4763 sw
tri 3242 4761 3244 4763 ne
rect 3244 4761 3683 4763
tri 3244 4710 3295 4761 ne
rect 3295 4731 3683 4761
rect 3919 4870 3968 4967
tri 3968 4870 4394 5296 sw
tri 4421 4870 4847 5296 ne
rect 4847 4910 5338 5296
tri 5338 4910 5724 5296 sw
tri 5791 4910 6177 5296 ne
rect 6177 5192 6711 5296
tri 6711 5192 6815 5296 sw
tri 7164 5192 7268 5296 ne
rect 7268 5241 7950 5296
rect 7268 5192 7589 5241
rect 6177 4910 6815 5192
tri 6815 4910 7097 5192 sw
tri 7268 4910 7550 5192 ne
rect 7550 5005 7589 5192
rect 7825 5188 7950 5241
rect 8186 5377 8266 5424
tri 8266 5377 8337 5448 sw
tri 8719 5377 8790 5448 ne
rect 8790 5377 11214 5448
rect 8186 5308 8337 5377
tri 8337 5308 8406 5377 sw
tri 8790 5308 8859 5377 ne
rect 8859 5364 11214 5377
tri 11214 5364 11347 5497 sw
rect 8859 5308 11347 5364
rect 8186 5192 8406 5308
tri 8406 5192 8522 5308 sw
tri 8859 5192 8975 5308 ne
rect 8975 5192 11347 5308
rect 8186 5188 8522 5192
rect 7825 5005 8522 5188
rect 7550 4910 8522 5005
rect 4847 4870 5724 4910
rect 3919 4846 4394 4870
rect 3919 4731 4131 4846
rect 3295 4710 4131 4731
rect 2757 4503 2842 4710
rect 1903 4466 2842 4503
rect 1903 4390 2139 4466
rect 0 4357 1449 4390
tri 1449 4357 1482 4390 sw
tri 1903 4357 1936 4390 ne
rect 1936 4357 2139 4390
rect 0 4333 1482 4357
rect 0 4097 294 4333
rect 530 4097 747 4333
rect 983 4097 1200 4333
rect 1436 4256 1482 4333
tri 1482 4256 1583 4357 sw
tri 1936 4256 2037 4357 ne
rect 2037 4256 2139 4357
rect 1436 4194 1583 4256
tri 1583 4194 1645 4256 sw
tri 2037 4194 2099 4256 ne
rect 2099 4230 2139 4256
rect 2375 4446 2842 4466
tri 2842 4446 3106 4710 sw
tri 3295 4446 3559 4710 ne
rect 3559 4639 4131 4710
rect 3559 4446 3683 4639
rect 2375 4417 3106 4446
tri 3106 4417 3135 4446 sw
tri 3559 4417 3588 4446 ne
rect 3588 4417 3683 4446
rect 2375 4412 3135 4417
rect 2375 4230 2521 4412
rect 2099 4194 2521 4230
rect 1436 4097 1645 4194
rect 0 4005 1645 4097
rect 0 3769 294 4005
rect 530 3769 747 4005
rect 983 3769 1200 4005
rect 1436 3769 1645 4005
rect 0 3740 1645 3769
tri 1645 3740 2099 4194 sw
tri 2099 3824 2469 4194 ne
rect 2469 4176 2521 4194
rect 2757 4393 3135 4412
rect 2757 4176 2867 4393
rect 2469 4157 2867 4176
rect 3103 4157 3135 4393
rect 2469 4084 3135 4157
rect 2469 3848 2521 4084
rect 2757 4066 3135 4084
rect 2757 3848 2867 4066
rect 2469 3830 2867 3848
rect 3103 4035 3135 4066
tri 3135 4035 3517 4417 sw
tri 3588 4379 3626 4417 ne
rect 3626 4403 3683 4417
rect 3919 4610 4131 4639
rect 4367 4843 4394 4846
tri 4394 4843 4421 4870 sw
tri 4847 4843 4874 4870 ne
rect 4874 4843 5724 4870
rect 4367 4710 4421 4843
tri 4421 4710 4554 4843 sw
tri 4874 4710 5007 4843 ne
rect 5007 4710 5724 4843
rect 4367 4610 4554 4710
rect 3919 4519 4554 4610
rect 3919 4403 4131 4519
rect 3626 4379 4131 4403
tri 3626 4035 3970 4379 ne
rect 3970 4283 4131 4379
rect 4367 4488 4554 4519
tri 4554 4488 4776 4710 sw
tri 5007 4488 5229 4710 ne
rect 5229 4488 5724 4710
rect 4367 4464 4776 4488
rect 4367 4283 4513 4464
rect 3970 4228 4513 4283
rect 4749 4446 4776 4464
tri 4776 4446 4818 4488 sw
tri 5229 4446 5271 4488 ne
rect 5271 4457 5724 4488
tri 5724 4457 6177 4910 sw
tri 6177 4457 6630 4910 ne
rect 6630 4855 7097 4910
tri 7097 4855 7152 4910 sw
tri 7550 4855 7605 4910 ne
rect 7605 4877 8522 4910
rect 7605 4855 7950 4877
rect 6630 4832 7152 4855
tri 7152 4832 7175 4855 sw
tri 7605 4832 7628 4855 ne
rect 7628 4832 7950 4855
rect 6630 4457 7175 4832
rect 5271 4446 6177 4457
rect 4749 4379 4818 4446
tri 4818 4379 4885 4446 sw
tri 5271 4379 5338 4446 ne
rect 5338 4379 6177 4446
tri 6177 4379 6255 4457 sw
tri 6630 4379 6708 4457 ne
rect 6708 4379 7175 4457
tri 7175 4379 7628 4832 sw
tri 7628 4617 7843 4832 ne
rect 7843 4641 7950 4832
rect 8186 4739 8522 4877
tri 8522 4739 8975 5192 sw
tri 8975 4739 9428 5192 ne
rect 9428 4739 11347 5192
rect 8186 4641 8975 4739
rect 7843 4620 8975 4641
tri 8975 4620 9094 4739 sw
tri 9428 4620 9547 4739 ne
rect 7843 4617 9094 4620
tri 7843 4379 8081 4617 ne
rect 8081 4487 9094 4617
tri 9094 4487 9227 4620 sw
rect 8081 4455 9227 4487
rect 8081 4379 8366 4455
rect 4749 4228 4885 4379
rect 3970 4191 4885 4228
rect 3970 4035 4131 4191
rect 3103 4011 3517 4035
rect 3103 3830 3249 4011
rect 2469 3824 3249 3830
tri 2469 3740 2553 3824 ne
rect 2553 3775 3249 3824
rect 3485 3993 3517 4011
tri 3517 3993 3559 4035 sw
tri 3970 3993 4012 4035 ne
rect 4012 3993 4131 4035
rect 3485 3775 3559 3993
rect 2553 3740 3559 3775
tri 1178 3420 1498 3740 ne
rect 1498 3451 2099 3740
tri 2099 3451 2388 3740 sw
tri 2553 3451 2842 3740 ne
rect 2842 3738 3559 3740
rect 2842 3502 2867 3738
rect 3103 3684 3559 3738
rect 3103 3502 3249 3684
rect 2842 3451 3249 3502
rect 1498 3420 2388 3451
rect 0 3362 1045 3420
rect 0 3126 757 3362
rect 993 3287 1045 3362
tri 1045 3287 1178 3420 sw
tri 1498 3287 1631 3420 ne
rect 1631 3287 2388 3420
rect 993 3272 1178 3287
tri 1178 3272 1193 3287 sw
tri 1631 3272 1646 3287 ne
rect 1646 3272 2388 3287
rect 993 3126 1193 3272
rect 0 2992 1193 3126
tri 1193 2992 1473 3272 sw
tri 1646 2992 1926 3272 ne
rect 1926 2997 2388 3272
tri 2388 2997 2842 3451 sw
tri 2842 3096 3197 3451 ne
rect 3197 3448 3249 3451
rect 3485 3656 3559 3684
tri 3559 3656 3896 3993 sw
tri 4012 3931 4074 3993 ne
rect 4074 3955 4131 3993
rect 4367 4137 4885 4191
rect 4367 3955 4513 4137
rect 4074 3931 4513 3955
tri 4074 3656 4349 3931 ne
rect 4349 3901 4513 3931
rect 4749 4090 4885 4137
tri 4885 4090 5174 4379 sw
tri 5338 4090 5627 4379 ne
rect 5627 4090 6255 4379
rect 4749 4066 5174 4090
rect 4749 3901 4911 4066
rect 4349 3830 4911 3901
rect 5147 3926 5174 4066
tri 5174 3926 5338 4090 sw
tri 5627 3926 5791 4090 ne
rect 5791 3990 6255 4090
tri 6255 3990 6644 4379 sw
tri 6708 3990 7097 4379 ne
rect 7097 4123 7628 4379
tri 7628 4123 7884 4379 sw
tri 8081 4123 8337 4379 ne
rect 8337 4219 8366 4379
rect 8602 4219 8956 4455
rect 9192 4219 9227 4455
rect 8337 4134 9227 4219
rect 7097 3990 7884 4123
tri 7884 3990 8017 4123 sw
rect 5791 3926 6644 3990
rect 5147 3830 5338 3926
rect 4349 3809 5338 3830
rect 4349 3656 4513 3809
rect 3485 3632 3896 3656
rect 3485 3448 3628 3632
rect 3197 3396 3628 3448
rect 3864 3575 3896 3632
tri 3896 3575 3977 3656 sw
tri 4349 3575 4430 3656 ne
rect 4430 3575 4513 3656
rect 3864 3451 3977 3575
tri 3977 3451 4101 3575 sw
tri 4430 3549 4456 3575 ne
rect 4456 3573 4513 3575
rect 4749 3739 5338 3809
rect 4749 3573 4911 3739
rect 4456 3549 4911 3573
tri 4456 3451 4554 3549 ne
rect 4554 3503 4911 3549
rect 5147 3575 5338 3739
tri 5338 3575 5689 3926 sw
tri 5791 3575 6142 3926 ne
rect 6142 3587 6644 3926
tri 6644 3587 7047 3990 sw
tri 7097 3720 7367 3990 ne
rect 7367 3962 8017 3990
rect 7367 3726 7402 3962
rect 7638 3726 7750 3962
rect 7986 3726 8017 3962
rect 6142 3575 7047 3587
rect 5147 3503 5689 3575
rect 4554 3462 5689 3503
tri 5689 3462 5802 3575 sw
tri 6142 3462 6255 3575 ne
rect 6255 3556 7047 3575
rect 6255 3462 6428 3556
rect 4554 3451 5802 3462
tri 5802 3451 5813 3462 sw
tri 6255 3451 6266 3462 ne
rect 6266 3451 6428 3462
rect 3864 3396 4101 3451
rect 3197 3356 4101 3396
rect 3197 3120 3249 3356
rect 3485 3305 4101 3356
rect 3485 3120 3628 3305
rect 3197 3096 3628 3120
tri 3197 2997 3296 3096 ne
rect 3296 3069 3628 3096
rect 3864 3187 4101 3305
tri 4101 3187 4365 3451 sw
tri 4554 3187 4818 3451 ne
rect 4818 3411 5813 3451
rect 4818 3187 4911 3411
rect 3864 3069 4365 3187
rect 3296 2997 4365 3069
rect 1926 2992 2842 2997
rect 0 2968 1473 2992
rect 0 2749 1151 2968
rect 0 2530 757 2749
tri 676 2489 717 2530 ne
rect 717 2513 757 2530
rect 993 2732 1151 2749
rect 1387 2819 1473 2968
tri 1473 2819 1646 2992 sw
tri 1926 2819 2099 2992 ne
rect 2099 2832 2842 2992
tri 2842 2832 3007 2997 sw
tri 3296 2832 3461 2997 ne
rect 3461 2977 4365 2997
rect 3461 2832 3628 2977
rect 2099 2819 3007 2832
tri 3007 2819 3020 2832 sw
tri 3461 2819 3474 2832 ne
rect 3474 2819 3628 2832
rect 1387 2732 1646 2819
rect 993 2668 1646 2732
tri 1646 2668 1797 2819 sw
tri 2099 2668 2250 2819 ne
rect 2250 2770 3020 2819
tri 3020 2770 3069 2819 sw
tri 3474 2770 3523 2819 ne
rect 3523 2770 3628 2819
rect 2250 2668 3069 2770
rect 993 2623 1797 2668
rect 993 2513 1496 2623
rect 717 2489 1496 2513
tri 717 2210 996 2489 ne
rect 996 2387 1496 2489
rect 1732 2530 1797 2623
tri 1797 2530 1935 2668 sw
tri 2250 2530 2388 2668 ne
rect 2388 2530 3069 2668
rect 1732 2387 1935 2530
rect 996 2366 1935 2387
tri 1935 2366 2099 2530 sw
tri 2388 2366 2552 2530 ne
rect 2552 2366 3069 2530
rect 996 2364 2099 2366
tri 2099 2364 2101 2366 sw
tri 2552 2364 2554 2366 ne
rect 2554 2364 3069 2366
rect 996 2355 2101 2364
rect 996 2210 1151 2355
rect 0 2076 542 2210
tri 542 2076 676 2210 sw
tri 996 2095 1111 2210 ne
rect 1111 2119 1151 2210
rect 1387 2119 2101 2355
rect 1111 2095 2101 2119
tri 1111 2076 1130 2095 ne
rect 1130 2076 2101 2095
rect 0 1863 676 2076
tri 676 1863 889 2076 sw
tri 1130 1863 1343 2076 ne
rect 1343 2010 2101 2076
rect 1343 1863 1496 2010
rect 0 1409 889 1863
tri 889 1409 1343 1863 sw
tri 1343 1750 1456 1863 ne
rect 1456 1774 1496 1863
rect 1732 1911 2101 2010
tri 2101 1911 2554 2364 sw
tri 2554 2316 2602 2364 ne
rect 2602 2316 3069 2364
tri 3069 2316 3523 2770 sw
tri 3523 2717 3576 2770 ne
rect 3576 2741 3628 2770
rect 3864 2818 4365 2977
tri 4365 2818 4734 3187 sw
tri 4818 3151 4854 3187 ne
rect 4854 3175 4911 3187
rect 5147 3187 5813 3411
tri 5813 3187 6077 3451 sw
tri 6266 3320 6397 3451 ne
rect 6397 3320 6428 3451
rect 6664 3320 6782 3556
rect 7018 3320 7047 3556
rect 5147 3175 6077 3187
rect 4854 3151 6077 3175
tri 4854 2818 5187 3151 ne
rect 5187 3146 6077 3151
rect 5187 2910 5233 3146
rect 5469 2910 5787 3146
rect 6023 2910 6077 3146
rect 3864 2741 4734 2818
rect 3576 2717 4734 2741
tri 3576 2316 3977 2717 ne
rect 3977 2685 4734 2717
tri 4734 2685 4867 2818 sw
rect 3977 2631 4867 2685
rect 3977 2395 4011 2631
rect 4247 2395 4597 2631
rect 4833 2395 4867 2631
tri 2602 1911 3007 2316 ne
rect 3007 2182 3523 2316
tri 3523 2182 3657 2316 sw
rect 3007 2129 3657 2182
rect 1732 1778 2554 1911
tri 2554 1778 2687 1911 sw
rect 1732 1774 2687 1778
rect 1456 1750 2687 1774
tri 1456 1409 1797 1750 ne
rect 1797 1721 2687 1750
rect 1797 1485 1836 1721
rect 2072 1485 2416 1721
rect 2652 1485 2687 1721
rect 0 1275 1343 1409
tri 1343 1275 1477 1409 sw
rect 0 1225 1477 1275
rect 0 1160 470 1225
tri 0 733 427 1160 ne
rect 427 989 470 1160
rect 706 989 834 1225
rect 1070 989 1198 1225
rect 1434 989 1477 1225
rect 427 749 1477 989
rect 427 513 470 749
rect 706 513 834 749
rect 1070 513 1198 749
rect 1434 513 1477 749
rect 427 272 1477 513
rect 427 36 470 272
rect 706 36 834 272
rect 1070 36 1198 272
rect 1434 36 1477 272
rect 427 0 1477 36
rect 1797 1358 2687 1485
rect 1797 1122 1836 1358
rect 2072 1122 2416 1358
rect 2652 1122 2687 1358
rect 1797 995 2687 1122
rect 1797 759 1836 995
rect 2072 759 2416 995
rect 2652 759 2687 995
rect 1797 631 2687 759
rect 1797 395 1836 631
rect 2072 395 2416 631
rect 2652 395 2687 631
rect 1797 267 2687 395
rect 1797 31 1836 267
rect 2072 31 2416 267
rect 2652 31 2687 267
rect 1797 0 2687 31
rect 3007 1893 3037 2129
rect 3273 1893 3393 2129
rect 3629 1893 3657 2129
rect 3007 1758 3657 1893
rect 3007 1522 3037 1758
rect 3273 1522 3393 1758
rect 3629 1522 3657 1758
rect 3007 1387 3657 1522
rect 3007 1151 3037 1387
rect 3273 1151 3393 1387
rect 3629 1151 3657 1387
rect 3007 1015 3657 1151
rect 3007 779 3037 1015
rect 3273 779 3393 1015
rect 3629 779 3657 1015
rect 3007 643 3657 779
rect 3007 407 3037 643
rect 3273 407 3393 643
rect 3629 407 3657 643
rect 3007 271 3657 407
rect 3007 35 3037 271
rect 3273 35 3393 271
rect 3629 35 3657 271
rect 3007 0 3657 35
rect 3977 2295 4867 2395
rect 3977 2059 4011 2295
rect 4247 2059 4597 2295
rect 4833 2059 4867 2295
rect 3977 1959 4867 2059
rect 3977 1723 4011 1959
rect 4247 1723 4597 1959
rect 4833 1723 4867 1959
rect 3977 1623 4867 1723
rect 3977 1387 4011 1623
rect 4247 1387 4597 1623
rect 4833 1387 4867 1623
rect 3977 1287 4867 1387
rect 3977 1051 4011 1287
rect 4247 1051 4597 1287
rect 4833 1051 4867 1287
rect 3977 951 4867 1051
rect 3977 715 4011 951
rect 4247 715 4597 951
rect 4833 715 4867 951
rect 3977 615 4867 715
rect 3977 379 4011 615
rect 4247 379 4597 615
rect 4833 379 4867 615
rect 3977 279 4867 379
rect 3977 43 4011 279
rect 4247 43 4597 279
rect 4833 43 4867 279
rect 3977 0 4867 43
rect 5187 2787 6077 2910
rect 5187 2551 5233 2787
rect 5469 2551 5787 2787
rect 6023 2551 6077 2787
rect 5187 2428 6077 2551
rect 5187 2192 5233 2428
rect 5469 2192 5787 2428
rect 6023 2192 6077 2428
rect 5187 2069 6077 2192
rect 5187 1833 5233 2069
rect 5469 1833 5787 2069
rect 6023 1833 6077 2069
rect 5187 1710 6077 1833
rect 5187 1474 5233 1710
rect 5469 1474 5787 1710
rect 6023 1474 6077 1710
rect 5187 1350 6077 1474
rect 5187 1114 5233 1350
rect 5469 1114 5787 1350
rect 6023 1114 6077 1350
rect 5187 990 6077 1114
rect 5187 754 5233 990
rect 5469 754 5787 990
rect 6023 754 6077 990
rect 5187 630 6077 754
rect 5187 394 5233 630
rect 5469 394 5787 630
rect 6023 394 6077 630
rect 5187 270 6077 394
rect 5187 34 5233 270
rect 5469 34 5787 270
rect 6023 34 6077 270
rect 5187 0 6077 34
rect 6397 3228 7047 3320
rect 6397 2992 6428 3228
rect 6664 2992 6782 3228
rect 7018 2992 7047 3228
rect 6397 2900 7047 2992
rect 6397 2664 6428 2900
rect 6664 2664 6782 2900
rect 7018 2664 7047 2900
rect 6397 2572 7047 2664
rect 6397 2336 6428 2572
rect 6664 2336 6782 2572
rect 7018 2336 7047 2572
rect 6397 2244 7047 2336
rect 6397 2008 6428 2244
rect 6664 2008 6782 2244
rect 7018 2008 7047 2244
rect 6397 1916 7047 2008
rect 6397 1680 6428 1916
rect 6664 1680 6782 1916
rect 7018 1680 7047 1916
rect 6397 1588 7047 1680
rect 6397 1352 6428 1588
rect 6664 1352 6782 1588
rect 7018 1352 7047 1588
rect 6397 1260 7047 1352
rect 6397 1024 6428 1260
rect 6664 1024 6782 1260
rect 7018 1024 7047 1260
rect 6397 931 7047 1024
rect 6397 695 6428 931
rect 6664 695 6782 931
rect 7018 695 7047 931
rect 6397 602 7047 695
rect 6397 366 6428 602
rect 6664 366 6782 602
rect 7018 366 7047 602
rect 6397 273 7047 366
rect 6397 37 6428 273
rect 6664 37 6782 273
rect 7018 37 7047 273
rect 6397 0 7047 37
rect 7367 3633 8017 3726
rect 7367 3397 7402 3633
rect 7638 3397 7750 3633
rect 7986 3397 8017 3633
rect 7367 3304 8017 3397
rect 7367 3068 7402 3304
rect 7638 3068 7750 3304
rect 7986 3068 8017 3304
rect 7367 2975 8017 3068
rect 7367 2739 7402 2975
rect 7638 2739 7750 2975
rect 7986 2739 8017 2975
rect 7367 2646 8017 2739
rect 7367 2410 7402 2646
rect 7638 2410 7750 2646
rect 7986 2410 8017 2646
rect 7367 2317 8017 2410
rect 7367 2081 7402 2317
rect 7638 2081 7750 2317
rect 7986 2081 8017 2317
rect 7367 1988 8017 2081
rect 7367 1752 7402 1988
rect 7638 1752 7750 1988
rect 7986 1752 8017 1988
rect 7367 1659 8017 1752
rect 7367 1423 7402 1659
rect 7638 1423 7750 1659
rect 7986 1423 8017 1659
rect 7367 1329 8017 1423
rect 7367 1093 7402 1329
rect 7638 1093 7750 1329
rect 7986 1093 8017 1329
rect 7367 999 8017 1093
rect 7367 763 7402 999
rect 7638 763 7750 999
rect 7986 763 8017 999
rect 7367 669 8017 763
rect 7367 433 7402 669
rect 7638 433 7750 669
rect 7986 433 8017 669
rect 7367 339 8017 433
rect 7367 103 7402 339
rect 7638 103 7750 339
rect 7986 103 8017 339
rect 7367 0 8017 103
rect 8337 3898 8366 4134
rect 8602 3898 8956 4134
rect 9192 3898 9227 4134
rect 8337 3813 9227 3898
rect 8337 3577 8366 3813
rect 8602 3577 8956 3813
rect 9192 3577 9227 3813
rect 8337 3492 9227 3577
rect 8337 3256 8366 3492
rect 8602 3256 8956 3492
rect 9192 3256 9227 3492
rect 8337 3171 9227 3256
rect 8337 2935 8366 3171
rect 8602 2935 8956 3171
rect 9192 2935 9227 3171
rect 8337 2849 9227 2935
rect 8337 2613 8366 2849
rect 8602 2613 8956 2849
rect 9192 2613 9227 2849
rect 8337 2527 9227 2613
rect 8337 2291 8366 2527
rect 8602 2291 8956 2527
rect 9192 2291 9227 2527
rect 8337 2205 9227 2291
rect 8337 1969 8366 2205
rect 8602 1969 8956 2205
rect 9192 1969 9227 2205
rect 8337 1883 9227 1969
rect 8337 1647 8366 1883
rect 8602 1647 8956 1883
rect 9192 1647 9227 1883
rect 8337 1561 9227 1647
rect 8337 1325 8366 1561
rect 8602 1325 8956 1561
rect 9192 1325 9227 1561
rect 8337 1239 9227 1325
rect 8337 1003 8366 1239
rect 8602 1003 8956 1239
rect 9192 1003 9227 1239
rect 8337 917 9227 1003
rect 8337 681 8366 917
rect 8602 681 8956 917
rect 9192 681 9227 917
rect 8337 595 9227 681
rect 8337 359 8366 595
rect 8602 359 8956 595
rect 9192 359 9227 595
rect 8337 273 9227 359
rect 8337 37 8366 273
rect 8602 37 8956 273
rect 9192 37 9227 273
rect 8337 0 9227 37
rect 9547 0 11347 4739
rect 11667 5487 12517 5576
rect 11667 5251 11703 5487
rect 11939 5251 12237 5487
rect 12473 5251 12517 5487
rect 11667 5162 12517 5251
rect 11667 4926 11703 5162
rect 11939 4926 12237 5162
rect 12473 4926 12517 5162
rect 11667 4837 12517 4926
rect 11667 4601 11703 4837
rect 11939 4601 12237 4837
rect 12473 4601 12517 4837
rect 11667 4512 12517 4601
rect 11667 4276 11703 4512
rect 11939 4276 12237 4512
rect 12473 4276 12517 4512
rect 11667 4187 12517 4276
rect 11667 3951 11703 4187
rect 11939 3951 12237 4187
rect 12473 3951 12517 4187
rect 11667 3862 12517 3951
rect 11667 3626 11703 3862
rect 11939 3626 12237 3862
rect 12473 3626 12517 3862
rect 11667 3537 12517 3626
rect 11667 3301 11703 3537
rect 11939 3301 12237 3537
rect 12473 3301 12517 3537
rect 11667 3211 12517 3301
rect 11667 2975 11703 3211
rect 11939 2975 12237 3211
rect 12473 2975 12517 3211
rect 11667 2885 12517 2975
rect 11667 2649 11703 2885
rect 11939 2649 12237 2885
rect 12473 2649 12517 2885
rect 11667 2559 12517 2649
rect 11667 2323 11703 2559
rect 11939 2323 12237 2559
rect 12473 2323 12517 2559
rect 11667 2233 12517 2323
rect 11667 1997 11703 2233
rect 11939 1997 12237 2233
rect 12473 1997 12517 2233
rect 11667 1907 12517 1997
rect 11667 1671 11703 1907
rect 11939 1671 12237 1907
rect 12473 1671 12517 1907
rect 11667 1581 12517 1671
rect 11667 1345 11703 1581
rect 11939 1345 12237 1581
rect 12473 1345 12517 1581
rect 11667 1255 12517 1345
rect 11667 1019 11703 1255
rect 11939 1019 12237 1255
rect 12473 1019 12517 1255
rect 11667 929 12517 1019
rect 11667 693 11703 929
rect 11939 693 12237 929
rect 12473 693 12517 929
rect 11667 603 12517 693
rect 11667 367 11703 603
rect 11939 367 12237 603
rect 12473 367 12517 603
rect 11667 277 12517 367
rect 11667 41 11703 277
rect 11939 41 12237 277
rect 12473 41 12517 277
rect 11667 0 12517 41
rect 12837 5948 13687 6043
rect 12837 5712 12869 5948
rect 13105 5712 13421 5948
rect 13657 5712 13687 5948
rect 12837 5617 13687 5712
rect 12837 5381 12869 5617
rect 13105 5381 13421 5617
rect 13657 5381 13687 5617
rect 12837 5286 13687 5381
rect 12837 5050 12869 5286
rect 13105 5050 13421 5286
rect 13657 5050 13687 5286
rect 12837 4955 13687 5050
rect 12837 4719 12869 4955
rect 13105 4719 13421 4955
rect 13657 4719 13687 4955
rect 12837 4624 13687 4719
rect 12837 4388 12869 4624
rect 13105 4388 13421 4624
rect 13657 4388 13687 4624
rect 12837 4293 13687 4388
rect 12837 4057 12869 4293
rect 13105 4057 13421 4293
rect 13657 4057 13687 4293
rect 12837 3962 13687 4057
rect 12837 3726 12869 3962
rect 13105 3726 13421 3962
rect 13657 3726 13687 3962
rect 12837 3631 13687 3726
rect 12837 3395 12869 3631
rect 13105 3395 13421 3631
rect 13657 3395 13687 3631
rect 12837 3300 13687 3395
rect 12837 3064 12869 3300
rect 13105 3064 13421 3300
rect 13657 3064 13687 3300
rect 12837 2969 13687 3064
rect 12837 2733 12869 2969
rect 13105 2733 13421 2969
rect 13657 2733 13687 2969
rect 12837 2638 13687 2733
rect 12837 2402 12869 2638
rect 13105 2402 13421 2638
rect 13657 2402 13687 2638
rect 12837 2307 13687 2402
rect 12837 2071 12869 2307
rect 13105 2071 13421 2307
rect 13657 2071 13687 2307
rect 12837 1976 13687 2071
rect 12837 1740 12869 1976
rect 13105 1740 13421 1976
rect 13657 1740 13687 1976
rect 12837 1644 13687 1740
rect 12837 1408 12869 1644
rect 13105 1408 13421 1644
rect 13657 1408 13687 1644
rect 12837 1312 13687 1408
rect 12837 1076 12869 1312
rect 13105 1076 13421 1312
rect 13657 1076 13687 1312
rect 12837 980 13687 1076
rect 12837 744 12869 980
rect 13105 744 13421 980
rect 13657 744 13687 980
rect 12837 648 13687 744
rect 12837 412 12869 648
rect 13105 412 13421 648
rect 13657 412 13687 648
rect 12837 316 13687 412
rect 12837 80 12869 316
rect 13105 80 13421 316
rect 13657 80 13687 316
rect 12837 0 13687 80
rect 14007 6253 14300 6489
rect 14536 6253 14624 6489
rect 14860 6253 14948 6489
rect 15184 6253 15272 6489
rect 15508 6253 15596 6489
rect 15832 6253 15920 6489
rect 16156 6253 16244 6489
rect 16480 6253 16568 6489
rect 16804 6253 16892 6489
rect 17128 6253 17216 6489
rect 17452 6253 17540 6489
rect 17776 6253 17864 6489
rect 18100 6253 18188 6489
rect 18424 6253 18512 6489
rect 18748 6253 18997 6489
rect 14007 6159 18997 6253
rect 14007 5923 14300 6159
rect 14536 5923 14624 6159
rect 14860 5923 14948 6159
rect 15184 5923 15272 6159
rect 15508 5923 15596 6159
rect 15832 5923 15920 6159
rect 16156 5923 16244 6159
rect 16480 5923 16568 6159
rect 16804 5923 16892 6159
rect 17128 5923 17216 6159
rect 17452 5923 17540 6159
rect 17776 5923 17864 6159
rect 18100 5923 18188 6159
rect 18424 5923 18512 6159
rect 18748 5923 18997 6159
rect 14007 5829 18997 5923
rect 14007 5593 14300 5829
rect 14536 5593 14624 5829
rect 14860 5593 14948 5829
rect 15184 5593 15272 5829
rect 15508 5593 15596 5829
rect 15832 5593 15920 5829
rect 16156 5593 16244 5829
rect 16480 5593 16568 5829
rect 16804 5593 16892 5829
rect 17128 5593 17216 5829
rect 17452 5593 17540 5829
rect 17776 5593 17864 5829
rect 18100 5593 18188 5829
rect 18424 5593 18512 5829
rect 18748 5593 18997 5829
rect 14007 5499 18997 5593
rect 14007 5263 14300 5499
rect 14536 5263 14624 5499
rect 14860 5263 14948 5499
rect 15184 5263 15272 5499
rect 15508 5263 15596 5499
rect 15832 5263 15920 5499
rect 16156 5263 16244 5499
rect 16480 5263 16568 5499
rect 16804 5263 16892 5499
rect 17128 5263 17216 5499
rect 17452 5263 17540 5499
rect 17776 5263 17864 5499
rect 18100 5263 18188 5499
rect 18424 5263 18512 5499
rect 18748 5263 18997 5499
rect 14007 5169 18997 5263
rect 14007 4933 14300 5169
rect 14536 4933 14624 5169
rect 14860 4933 14948 5169
rect 15184 4933 15272 5169
rect 15508 4933 15596 5169
rect 15832 4933 15920 5169
rect 16156 4933 16244 5169
rect 16480 4933 16568 5169
rect 16804 4933 16892 5169
rect 17128 4933 17216 5169
rect 17452 4933 17540 5169
rect 17776 4933 17864 5169
rect 18100 4933 18188 5169
rect 18424 4933 18512 5169
rect 18748 4933 18997 5169
rect 14007 4839 18997 4933
rect 14007 4603 14300 4839
rect 14536 4603 14624 4839
rect 14860 4603 14948 4839
rect 15184 4603 15272 4839
rect 15508 4603 15596 4839
rect 15832 4603 15920 4839
rect 16156 4603 16244 4839
rect 16480 4603 16568 4839
rect 16804 4603 16892 4839
rect 17128 4603 17216 4839
rect 17452 4603 17540 4839
rect 17776 4603 17864 4839
rect 18100 4603 18188 4839
rect 18424 4603 18512 4839
rect 18748 4603 18997 4839
rect 14007 4509 18997 4603
rect 14007 4273 14300 4509
rect 14536 4273 14624 4509
rect 14860 4273 14948 4509
rect 15184 4273 15272 4509
rect 15508 4273 15596 4509
rect 15832 4273 15920 4509
rect 16156 4273 16244 4509
rect 16480 4273 16568 4509
rect 16804 4273 16892 4509
rect 17128 4273 17216 4509
rect 17452 4273 17540 4509
rect 17776 4273 17864 4509
rect 18100 4273 18188 4509
rect 18424 4273 18512 4509
rect 18748 4273 18997 4509
rect 14007 4179 18997 4273
rect 14007 3943 14300 4179
rect 14536 3943 14624 4179
rect 14860 3943 14948 4179
rect 15184 3943 15272 4179
rect 15508 3943 15596 4179
rect 15832 3943 15920 4179
rect 16156 3943 16244 4179
rect 16480 3943 16568 4179
rect 16804 3943 16892 4179
rect 17128 3943 17216 4179
rect 17452 3943 17540 4179
rect 17776 3943 17864 4179
rect 18100 3943 18188 4179
rect 18424 3943 18512 4179
rect 18748 3943 18997 4179
rect 14007 3849 18997 3943
rect 14007 3613 14300 3849
rect 14536 3613 14624 3849
rect 14860 3613 14948 3849
rect 15184 3613 15272 3849
rect 15508 3613 15596 3849
rect 15832 3613 15920 3849
rect 16156 3613 16244 3849
rect 16480 3613 16568 3849
rect 16804 3613 16892 3849
rect 17128 3613 17216 3849
rect 17452 3613 17540 3849
rect 17776 3613 17864 3849
rect 18100 3613 18188 3849
rect 18424 3613 18512 3849
rect 18748 3613 18997 3849
rect 14007 3519 18997 3613
rect 14007 3283 14300 3519
rect 14536 3283 14624 3519
rect 14860 3283 14948 3519
rect 15184 3283 15272 3519
rect 15508 3283 15596 3519
rect 15832 3283 15920 3519
rect 16156 3283 16244 3519
rect 16480 3283 16568 3519
rect 16804 3283 16892 3519
rect 17128 3283 17216 3519
rect 17452 3283 17540 3519
rect 17776 3283 17864 3519
rect 18100 3283 18188 3519
rect 18424 3283 18512 3519
rect 18748 3283 18997 3519
rect 14007 3188 18997 3283
rect 14007 2952 14300 3188
rect 14536 2952 14624 3188
rect 14860 2952 14948 3188
rect 15184 2952 15272 3188
rect 15508 2952 15596 3188
rect 15832 2952 15920 3188
rect 16156 2952 16244 3188
rect 16480 2952 16568 3188
rect 16804 2952 16892 3188
rect 17128 2952 17216 3188
rect 17452 2952 17540 3188
rect 17776 2952 17864 3188
rect 18100 2952 18188 3188
rect 18424 2952 18512 3188
rect 18748 2952 18997 3188
rect 14007 2857 18997 2952
rect 14007 2621 14300 2857
rect 14536 2621 14624 2857
rect 14860 2621 14948 2857
rect 15184 2621 15272 2857
rect 15508 2621 15596 2857
rect 15832 2621 15920 2857
rect 16156 2621 16244 2857
rect 16480 2621 16568 2857
rect 16804 2621 16892 2857
rect 17128 2621 17216 2857
rect 17452 2621 17540 2857
rect 17776 2621 17864 2857
rect 18100 2621 18188 2857
rect 18424 2621 18512 2857
rect 18748 2621 18997 2857
rect 14007 2526 18997 2621
rect 14007 2290 14300 2526
rect 14536 2290 14624 2526
rect 14860 2290 14948 2526
rect 15184 2290 15272 2526
rect 15508 2290 15596 2526
rect 15832 2290 15920 2526
rect 16156 2290 16244 2526
rect 16480 2290 16568 2526
rect 16804 2290 16892 2526
rect 17128 2290 17216 2526
rect 17452 2290 17540 2526
rect 17776 2290 17864 2526
rect 18100 2290 18188 2526
rect 18424 2290 18512 2526
rect 18748 2290 18997 2526
rect 14007 2195 18997 2290
rect 14007 1959 14300 2195
rect 14536 1959 14624 2195
rect 14860 1959 14948 2195
rect 15184 1959 15272 2195
rect 15508 1959 15596 2195
rect 15832 1959 15920 2195
rect 16156 1959 16244 2195
rect 16480 1959 16568 2195
rect 16804 1959 16892 2195
rect 17128 1959 17216 2195
rect 17452 1959 17540 2195
rect 17776 1959 17864 2195
rect 18100 1959 18188 2195
rect 18424 1959 18512 2195
rect 18748 1959 18997 2195
rect 14007 1864 18997 1959
rect 14007 1628 14300 1864
rect 14536 1628 14624 1864
rect 14860 1628 14948 1864
rect 15184 1628 15272 1864
rect 15508 1628 15596 1864
rect 15832 1628 15920 1864
rect 16156 1628 16244 1864
rect 16480 1628 16568 1864
rect 16804 1628 16892 1864
rect 17128 1628 17216 1864
rect 17452 1628 17540 1864
rect 17776 1628 17864 1864
rect 18100 1628 18188 1864
rect 18424 1628 18512 1864
rect 18748 1628 18997 1864
rect 14007 1533 18997 1628
rect 14007 1297 14300 1533
rect 14536 1297 14624 1533
rect 14860 1297 14948 1533
rect 15184 1297 15272 1533
rect 15508 1297 15596 1533
rect 15832 1297 15920 1533
rect 16156 1297 16244 1533
rect 16480 1297 16568 1533
rect 16804 1297 16892 1533
rect 17128 1297 17216 1533
rect 17452 1297 17540 1533
rect 17776 1297 17864 1533
rect 18100 1297 18188 1533
rect 18424 1297 18512 1533
rect 18748 1297 18997 1533
rect 14007 1202 18997 1297
rect 14007 966 14300 1202
rect 14536 966 14624 1202
rect 14860 966 14948 1202
rect 15184 966 15272 1202
rect 15508 966 15596 1202
rect 15832 966 15920 1202
rect 16156 966 16244 1202
rect 16480 966 16568 1202
rect 16804 966 16892 1202
rect 17128 966 17216 1202
rect 17452 966 17540 1202
rect 17776 966 17864 1202
rect 18100 966 18188 1202
rect 18424 966 18512 1202
rect 18748 966 18997 1202
rect 14007 871 18997 966
rect 14007 635 14300 871
rect 14536 635 14624 871
rect 14860 635 14948 871
rect 15184 635 15272 871
rect 15508 635 15596 871
rect 15832 635 15920 871
rect 16156 635 16244 871
rect 16480 635 16568 871
rect 16804 635 16892 871
rect 17128 635 17216 871
rect 17452 635 17540 871
rect 17776 635 17864 871
rect 18100 635 18188 871
rect 18424 635 18512 871
rect 18748 635 18997 871
rect 14007 540 18997 635
rect 14007 304 14300 540
rect 14536 304 14624 540
rect 14860 304 14948 540
rect 15184 304 15272 540
rect 15508 304 15596 540
rect 15832 304 15920 540
rect 16156 304 16244 540
rect 16480 304 16568 540
rect 16804 304 16892 540
rect 17128 304 17216 540
rect 17452 304 17540 540
rect 17776 304 17864 540
rect 18100 304 18188 540
rect 18424 304 18512 540
rect 18748 304 18997 540
rect 14007 0 18997 304
rect 35157 8462 40000 8548
rect 35157 8226 35250 8462
rect 35486 8226 35584 8462
rect 35820 8226 35918 8462
rect 36154 8226 36252 8462
rect 36488 8226 36586 8462
rect 36822 8226 36920 8462
rect 37156 8226 37254 8462
rect 37490 8226 37588 8462
rect 37824 8226 37922 8462
rect 38158 8226 38256 8462
rect 38492 8226 38590 8462
rect 38826 8226 38924 8462
rect 39160 8226 39258 8462
rect 39494 8226 39592 8462
rect 39828 8226 40000 8462
rect 35157 8140 40000 8226
rect 35157 7904 35250 8140
rect 35486 7904 35584 8140
rect 35820 7904 35918 8140
rect 36154 7904 36252 8140
rect 36488 7904 36586 8140
rect 36822 7904 36920 8140
rect 37156 7904 37254 8140
rect 37490 7904 37588 8140
rect 37824 7904 37922 8140
rect 38158 7904 38256 8140
rect 38492 7904 38590 8140
rect 38826 7904 38924 8140
rect 39160 7904 39258 8140
rect 39494 7904 39592 8140
rect 39828 7904 40000 8140
rect 35157 7818 40000 7904
rect 35157 7582 35250 7818
rect 35486 7582 35584 7818
rect 35820 7582 35918 7818
rect 36154 7582 36252 7818
rect 36488 7582 36586 7818
rect 36822 7582 36920 7818
rect 37156 7582 37254 7818
rect 37490 7582 37588 7818
rect 37824 7582 37922 7818
rect 38158 7582 38256 7818
rect 38492 7582 38590 7818
rect 38826 7582 38924 7818
rect 39160 7582 39258 7818
rect 39494 7582 39592 7818
rect 39828 7582 40000 7818
rect 35157 7496 40000 7582
rect 35157 7260 35250 7496
rect 35486 7260 35584 7496
rect 35820 7260 35918 7496
rect 36154 7260 36252 7496
rect 36488 7260 36586 7496
rect 36822 7260 36920 7496
rect 37156 7260 37254 7496
rect 37490 7260 37588 7496
rect 37824 7260 37922 7496
rect 38158 7260 38256 7496
rect 38492 7260 38590 7496
rect 38826 7260 38924 7496
rect 39160 7260 39258 7496
rect 39494 7260 39592 7496
rect 39828 7260 40000 7496
rect 35157 7174 40000 7260
rect 35157 6938 35250 7174
rect 35486 6938 35584 7174
rect 35820 6938 35918 7174
rect 36154 6938 36252 7174
rect 36488 6938 36586 7174
rect 36822 6938 36920 7174
rect 37156 6938 37254 7174
rect 37490 6938 37588 7174
rect 37824 6938 37922 7174
rect 38158 6938 38256 7174
rect 38492 6938 38590 7174
rect 38826 6938 38924 7174
rect 39160 6938 39258 7174
rect 39494 6938 39592 7174
rect 39828 6938 40000 7174
rect 35157 6852 40000 6938
rect 35157 6616 35250 6852
rect 35486 6616 35584 6852
rect 35820 6616 35918 6852
rect 36154 6616 36252 6852
rect 36488 6616 36586 6852
rect 36822 6616 36920 6852
rect 37156 6616 37254 6852
rect 37490 6616 37588 6852
rect 37824 6616 37922 6852
rect 38158 6616 38256 6852
rect 38492 6616 38590 6852
rect 38826 6616 38924 6852
rect 39160 6616 39258 6852
rect 39494 6616 39592 6852
rect 39828 6616 40000 6852
rect 35157 6530 40000 6616
rect 35157 6294 35250 6530
rect 35486 6294 35584 6530
rect 35820 6294 35918 6530
rect 36154 6294 36252 6530
rect 36488 6294 36586 6530
rect 36822 6294 36920 6530
rect 37156 6294 37254 6530
rect 37490 6294 37588 6530
rect 37824 6294 37922 6530
rect 38158 6294 38256 6530
rect 38492 6294 38590 6530
rect 38826 6294 38924 6530
rect 39160 6294 39258 6530
rect 39494 6294 39592 6530
rect 39828 6294 40000 6530
rect 35157 6208 40000 6294
rect 35157 5972 35250 6208
rect 35486 5972 35584 6208
rect 35820 5972 35918 6208
rect 36154 5972 36252 6208
rect 36488 5972 36586 6208
rect 36822 5972 36920 6208
rect 37156 5972 37254 6208
rect 37490 5972 37588 6208
rect 37824 5972 37922 6208
rect 38158 5972 38256 6208
rect 38492 5972 38590 6208
rect 38826 5972 38924 6208
rect 39160 5972 39258 6208
rect 39494 5972 39592 6208
rect 39828 5972 40000 6208
rect 35157 5886 40000 5972
rect 35157 5650 35250 5886
rect 35486 5650 35584 5886
rect 35820 5650 35918 5886
rect 36154 5650 36252 5886
rect 36488 5650 36586 5886
rect 36822 5650 36920 5886
rect 37156 5650 37254 5886
rect 37490 5650 37588 5886
rect 37824 5650 37922 5886
rect 38158 5650 38256 5886
rect 38492 5650 38590 5886
rect 38826 5650 38924 5886
rect 39160 5650 39258 5886
rect 39494 5650 39592 5886
rect 39828 5650 40000 5886
rect 35157 5564 40000 5650
rect 35157 5328 35250 5564
rect 35486 5328 35584 5564
rect 35820 5328 35918 5564
rect 36154 5328 36252 5564
rect 36488 5328 36586 5564
rect 36822 5328 36920 5564
rect 37156 5328 37254 5564
rect 37490 5328 37588 5564
rect 37824 5328 37922 5564
rect 38158 5328 38256 5564
rect 38492 5328 38590 5564
rect 38826 5328 38924 5564
rect 39160 5328 39258 5564
rect 39494 5328 39592 5564
rect 39828 5328 40000 5564
rect 35157 5242 40000 5328
rect 35157 5006 35250 5242
rect 35486 5006 35584 5242
rect 35820 5006 35918 5242
rect 36154 5006 36252 5242
rect 36488 5006 36586 5242
rect 36822 5006 36920 5242
rect 37156 5006 37254 5242
rect 37490 5006 37588 5242
rect 37824 5006 37922 5242
rect 38158 5006 38256 5242
rect 38492 5006 38590 5242
rect 38826 5006 38924 5242
rect 39160 5006 39258 5242
rect 39494 5006 39592 5242
rect 39828 5006 40000 5242
rect 35157 4920 40000 5006
rect 35157 4684 35250 4920
rect 35486 4684 35584 4920
rect 35820 4684 35918 4920
rect 36154 4684 36252 4920
rect 36488 4684 36586 4920
rect 36822 4684 36920 4920
rect 37156 4684 37254 4920
rect 37490 4684 37588 4920
rect 37824 4684 37922 4920
rect 38158 4684 38256 4920
rect 38492 4684 38590 4920
rect 38826 4684 38924 4920
rect 39160 4684 39258 4920
rect 39494 4684 39592 4920
rect 39828 4684 40000 4920
rect 35157 4598 40000 4684
rect 35157 4362 35250 4598
rect 35486 4362 35584 4598
rect 35820 4362 35918 4598
rect 36154 4362 36252 4598
rect 36488 4362 36586 4598
rect 36822 4362 36920 4598
rect 37156 4362 37254 4598
rect 37490 4362 37588 4598
rect 37824 4362 37922 4598
rect 38158 4362 38256 4598
rect 38492 4362 38590 4598
rect 38826 4362 38924 4598
rect 39160 4362 39258 4598
rect 39494 4362 39592 4598
rect 39828 4362 40000 4598
rect 35157 4276 40000 4362
rect 35157 4040 35250 4276
rect 35486 4040 35584 4276
rect 35820 4040 35918 4276
rect 36154 4040 36252 4276
rect 36488 4040 36586 4276
rect 36822 4040 36920 4276
rect 37156 4040 37254 4276
rect 37490 4040 37588 4276
rect 37824 4040 37922 4276
rect 38158 4040 38256 4276
rect 38492 4040 38590 4276
rect 38826 4040 38924 4276
rect 39160 4040 39258 4276
rect 39494 4040 39592 4276
rect 39828 4040 40000 4276
rect 35157 3954 40000 4040
rect 35157 3718 35250 3954
rect 35486 3718 35584 3954
rect 35820 3718 35918 3954
rect 36154 3718 36252 3954
rect 36488 3718 36586 3954
rect 36822 3718 36920 3954
rect 37156 3718 37254 3954
rect 37490 3718 37588 3954
rect 37824 3718 37922 3954
rect 38158 3718 38256 3954
rect 38492 3718 38590 3954
rect 38826 3718 38924 3954
rect 39160 3718 39258 3954
rect 39494 3718 39592 3954
rect 39828 3718 40000 3954
rect 35157 3632 40000 3718
rect 35157 3396 35250 3632
rect 35486 3396 35584 3632
rect 35820 3396 35918 3632
rect 36154 3396 36252 3632
rect 36488 3396 36586 3632
rect 36822 3396 36920 3632
rect 37156 3396 37254 3632
rect 37490 3396 37588 3632
rect 37824 3396 37922 3632
rect 38158 3396 38256 3632
rect 38492 3396 38590 3632
rect 38826 3396 38924 3632
rect 39160 3396 39258 3632
rect 39494 3396 39592 3632
rect 39828 3396 40000 3632
rect 35157 3310 40000 3396
rect 35157 3074 35250 3310
rect 35486 3074 35584 3310
rect 35820 3074 35918 3310
rect 36154 3074 36252 3310
rect 36488 3074 36586 3310
rect 36822 3074 36920 3310
rect 37156 3074 37254 3310
rect 37490 3074 37588 3310
rect 37824 3074 37922 3310
rect 38158 3074 38256 3310
rect 38492 3074 38590 3310
rect 38826 3074 38924 3310
rect 39160 3074 39258 3310
rect 39494 3074 39592 3310
rect 39828 3074 40000 3310
rect 35157 2987 40000 3074
rect 35157 2751 35250 2987
rect 35486 2751 35584 2987
rect 35820 2751 35918 2987
rect 36154 2751 36252 2987
rect 36488 2751 36586 2987
rect 36822 2751 36920 2987
rect 37156 2751 37254 2987
rect 37490 2751 37588 2987
rect 37824 2751 37922 2987
rect 38158 2751 38256 2987
rect 38492 2751 38590 2987
rect 38826 2751 38924 2987
rect 39160 2751 39258 2987
rect 39494 2751 39592 2987
rect 39828 2751 40000 2987
rect 35157 2664 40000 2751
rect 35157 2428 35250 2664
rect 35486 2428 35584 2664
rect 35820 2428 35918 2664
rect 36154 2428 36252 2664
rect 36488 2428 36586 2664
rect 36822 2428 36920 2664
rect 37156 2428 37254 2664
rect 37490 2428 37588 2664
rect 37824 2428 37922 2664
rect 38158 2428 38256 2664
rect 38492 2428 38590 2664
rect 38826 2428 38924 2664
rect 39160 2428 39258 2664
rect 39494 2428 39592 2664
rect 39828 2428 40000 2664
rect 35157 2341 40000 2428
rect 35157 2105 35250 2341
rect 35486 2105 35584 2341
rect 35820 2105 35918 2341
rect 36154 2105 36252 2341
rect 36488 2105 36586 2341
rect 36822 2105 36920 2341
rect 37156 2105 37254 2341
rect 37490 2105 37588 2341
rect 37824 2105 37922 2341
rect 38158 2105 38256 2341
rect 38492 2105 38590 2341
rect 38826 2105 38924 2341
rect 39160 2105 39258 2341
rect 39494 2105 39592 2341
rect 39828 2105 40000 2341
rect 35157 2018 40000 2105
rect 35157 1782 35250 2018
rect 35486 1782 35584 2018
rect 35820 1782 35918 2018
rect 36154 1782 36252 2018
rect 36488 1782 36586 2018
rect 36822 1782 36920 2018
rect 37156 1782 37254 2018
rect 37490 1782 37588 2018
rect 37824 1782 37922 2018
rect 38158 1782 38256 2018
rect 38492 1782 38590 2018
rect 38826 1782 38924 2018
rect 39160 1782 39258 2018
rect 39494 1782 39592 2018
rect 39828 1782 40000 2018
rect 35157 1695 40000 1782
rect 35157 1459 35250 1695
rect 35486 1459 35584 1695
rect 35820 1459 35918 1695
rect 36154 1459 36252 1695
rect 36488 1459 36586 1695
rect 36822 1459 36920 1695
rect 37156 1459 37254 1695
rect 37490 1459 37588 1695
rect 37824 1459 37922 1695
rect 38158 1459 38256 1695
rect 38492 1459 38590 1695
rect 38826 1459 38924 1695
rect 39160 1459 39258 1695
rect 39494 1459 39592 1695
rect 39828 1459 40000 1695
rect 35157 1372 40000 1459
rect 35157 1136 35250 1372
rect 35486 1136 35584 1372
rect 35820 1136 35918 1372
rect 36154 1136 36252 1372
rect 36488 1136 36586 1372
rect 36822 1136 36920 1372
rect 37156 1136 37254 1372
rect 37490 1136 37588 1372
rect 37824 1136 37922 1372
rect 38158 1136 38256 1372
rect 38492 1136 38590 1372
rect 38826 1136 38924 1372
rect 39160 1136 39258 1372
rect 39494 1136 39592 1372
rect 39828 1136 40000 1372
rect 35157 1049 40000 1136
rect 35157 813 35250 1049
rect 35486 813 35584 1049
rect 35820 813 35918 1049
rect 36154 813 36252 1049
rect 36488 813 36586 1049
rect 36822 813 36920 1049
rect 37156 813 37254 1049
rect 37490 813 37588 1049
rect 37824 813 37922 1049
rect 38158 813 38256 1049
rect 38492 813 38590 1049
rect 38826 813 38924 1049
rect 39160 813 39258 1049
rect 39494 813 39592 1049
rect 39828 813 40000 1049
rect 35157 726 40000 813
rect 35157 490 35250 726
rect 35486 490 35584 726
rect 35820 490 35918 726
rect 36154 490 36252 726
rect 36488 490 36586 726
rect 36822 490 36920 726
rect 37156 490 37254 726
rect 37490 490 37588 726
rect 37824 490 37922 726
rect 38158 490 38256 726
rect 38492 490 38590 726
rect 38826 490 38924 726
rect 39160 490 39258 726
rect 39494 490 39592 726
rect 39828 490 40000 726
rect 35157 403 40000 490
rect 35157 167 35250 403
rect 35486 167 35584 403
rect 35820 167 35918 403
rect 36154 167 36252 403
rect 36488 167 36586 403
rect 36822 167 36920 403
rect 37156 167 37254 403
rect 37490 167 37588 403
rect 37824 167 37922 403
rect 38158 167 38256 403
rect 38492 167 38590 403
rect 38826 167 38924 403
rect 39160 167 39258 403
rect 39494 167 39592 403
rect 39828 167 40000 403
rect 35157 0 40000 167
<< labels >>
flabel metal5 s 0 10280 254 12080 3 FreeSans 520 0 0 0 VSSA
port 1 nsew signal bidirectional
flabel metal5 s 127 11138 127 11138 3 FreeSans 520 180 0 0 VSSA
flabel metal5 s 0 35890 254 40733 3 FreeSans 520 180 0 0 VSSIO
port 2 nsew signal bidirectional
flabel metal5 s 0 7130 254 7780 3 FreeSans 520 180 0 0 VSWITCH
port 3 nsew signal bidirectional
flabel metal5 s 0 5920 254 6810 3 FreeSans 520 180 0 0 VSSIO
port 2 nsew signal bidirectional
flabel metal5 s 0 9070 254 9960 3 FreeSans 520 180 0 0 VSSD
port 4 nsew signal bidirectional
flabel metal5 s 0 8101 254 8750 3 FreeSans 520 180 0 0 VSSA
port 1 nsew
flabel metal5 s 0 12400 254 13250 3 FreeSans 520 180 0 0 VSSIO_Q
port 5 nsew signal bidirectional
flabel metal5 s 0 13570 254 14420 3 FreeSans 520 180 0 0 VDDIO_Q
port 6 nsew signal bidirectional
flabel metal5 s 0 14740 254 19730 3 FreeSans 520 180 0 0 VDDIO
port 7 nsew signal bidirectional
flabel metal5 s 0 3740 251 4390 3 FreeSans 520 180 0 0 VDDA
port 8 nsew signal bidirectional
flabel metal5 s 0 1160 254 2210 3 FreeSans 520 180 0 0 VCCHIB
port 9 nsew signal bidirectional
flabel metal5 s 0 2530 254 3420 3 FreeSans 520 180 0 0 VCCD
port 10 nsew signal bidirectional
flabel metal5 s 0 4710 254 5600 3 FreeSans 520 180 0 0 VDDIO
port 7 nsew signal bidirectional
flabel metal5 s 3977 0 4867 254 3 FreeSans 520 270 0 0 VDDIO
port 7 nsew signal bidirectional
flabel metal5 s 1797 0 2687 254 3 FreeSans 520 270 0 0 VCCD
port 10 nsew signal bidirectional
flabel metal5 s 427 0 1477 254 3 FreeSans 520 270 0 0 VCCHIB
port 9 nsew signal bidirectional
flabel metal5 s 3007 0 3657 251 3 FreeSans 520 270 0 0 VDDA
port 8 nsew signal bidirectional
flabel metal5 s 14007 0 18997 254 3 FreeSans 520 270 0 0 VDDIO
port 7 nsew signal bidirectional
flabel metal5 s 12837 0 13687 254 3 FreeSans 520 270 0 0 VDDIO_Q
port 6 nsew signal bidirectional
flabel metal5 s 11667 0 12517 254 3 FreeSans 520 270 0 0 VSSIO_Q
port 5 nsew signal bidirectional
flabel metal5 s 7368 0 8017 254 3 FreeSans 520 270 0 0 VSSA
port 1 nsew
flabel metal5 s 8337 0 9227 254 3 FreeSans 520 270 0 0 VSSD
port 4 nsew signal bidirectional
flabel metal5 s 5187 0 6077 254 3 FreeSans 520 270 0 0 VSSIO
port 2 nsew signal bidirectional
flabel metal5 s 6397 0 7047 254 3 FreeSans 520 270 0 0 VSWITCH
port 3 nsew signal bidirectional
flabel metal5 s 35157 0 40000 254 3 FreeSans 520 270 0 0 VSSIO
port 2 nsew signal bidirectional
flabel metal5 s 9547 0 11347 254 3 FreeSans 520 270 0 0 VSSA
port 1 nsew
flabel metal5 s 10258 127 10258 127 3 FreeSans 520 90 0 0 VSSA
flabel metal4 s 0 11358 100 11954 3 FreeSans 520 0 0 0 AMUXBUS_A
port 11 nsew signal bidirectional
flabel metal4 s 0 10406 115 11002 3 FreeSans 520 0 0 0 AMUXBUS_B
port 12 nsew signal bidirectional
flabel metal4 s 0 10280 254 10346 3 FreeSans 520 0 0 0 VSSA
port 1 nsew
flabel metal4 s 0 1140 254 2230 3 FreeSans 520 180 0 0 VCCHIB
port 9 nsew signal bidirectional
flabel metal4 s 0 2510 254 3440 3 FreeSans 520 180 0 0 VCCD
port 10 nsew signal bidirectional
flabel metal4 s 0 3720 251 4410 3 FreeSans 520 180 0 0 VDDA
port 8 nsew signal bidirectional
flabel metal4 s 0 4690 254 5620 3 FreeSans 520 180 0 0 VDDIO
port 7 nsew signal bidirectional
flabel metal4 s 0 5900 254 6830 3 FreeSans 520 180 0 0 VSSIO
port 2 nsew signal bidirectional
flabel metal4 s 0 7110 254 7800 3 FreeSans 520 180 0 0 VSWITCH
port 3 nsew signal bidirectional
flabel metal4 s 0 8080 254 8770 3 FreeSans 520 180 0 0 VSSA
port 1 nsew
flabel metal4 s 0 9050 254 9980 3 FreeSans 520 180 0 0 VSSD
port 4 nsew signal bidirectional
flabel metal4 s 0 11062 254 11298 3 FreeSans 520 0 0 0 VSSA
port 1 nsew
flabel metal4 s 0 12014 254 12080 3 FreeSans 520 0 0 0 VSSA
port 1 nsew
flabel metal4 s 0 12380 254 13270 3 FreeSans 520 180 0 0 VSSIO_Q
port 5 nsew signal bidirectional
flabel metal4 s 0 13550 254 14440 3 FreeSans 520 180 0 0 VDDIO_Q
port 6 nsew signal bidirectional
flabel metal4 s 0 14741 254 19733 3 FreeSans 520 180 0 0 VDDIO
port 7 nsew signal bidirectional
flabel metal4 s 0 35890 254 40733 3 FreeSans 520 180 0 0 VSSIO
port 2 nsew signal bidirectional
flabel metal4 s 127 38907 127 38907 3 FreeSans 520 180 0 0 VSSIO
flabel metal4 s 35157 0 40000 254 3 FreeSans 520 270 0 0 VSSIO
port 2 nsew
flabel metal4 s 38174 127 38174 127 3 FreeSans 520 270 0 0 VSSIO
flabel metal4 s 14008 0 19000 254 3 FreeSans 520 270 0 0 VDDIO
port 7 nsew signal bidirectional
flabel metal4 s 12817 0 13707 254 3 FreeSans 520 270 0 0 VDDIO_Q
port 6 nsew signal bidirectional
flabel metal4 s 11647 0 12537 254 3 FreeSans 520 270 0 0 VSSIO_Q
port 5 nsew signal bidirectional
flabel metal4 s 11281 0 11347 254 3 FreeSans 520 90 0 0 VSSA
port 1 nsew
flabel metal4 s 10329 0 10565 254 3 FreeSans 520 90 0 0 VSSA
port 1 nsew
flabel metal4 s 8317 0 9247 254 3 FreeSans 520 270 0 0 VSSD
port 4 nsew signal bidirectional
flabel metal4 s 7347 0 8037 254 3 FreeSans 520 270 0 0 VSSA
port 1 nsew
flabel metal4 s 6377 0 7067 254 3 FreeSans 520 270 0 0 VSWITCH
port 3 nsew signal bidirectional
flabel metal4 s 5167 0 6097 254 3 FreeSans 520 270 0 0 VSSIO
port 2 nsew
flabel metal4 s 3957 0 4887 254 3 FreeSans 520 270 0 0 VDDIO
port 7 nsew signal bidirectional
flabel metal4 s 2987 0 3677 251 3 FreeSans 520 270 0 0 VDDA
port 8 nsew signal bidirectional
flabel metal4 s 1777 0 2707 254 3 FreeSans 520 270 0 0 VCCD
port 10 nsew signal bidirectional
flabel metal4 s 407 0 1497 254 3 FreeSans 520 270 0 0 VCCHIB
port 9 nsew signal bidirectional
flabel metal4 s 9547 0 9613 254 3 FreeSans 520 90 0 0 VSSA
port 1 nsew
flabel metal4 s 10625 0 11221 100 3 FreeSans 520 90 0 0 AMUXBUS_A
port 11 nsew signal bidirectional
flabel metal4 s 9673 0 10269 115 3 FreeSans 520 90 0 0 AMUXBUS_B
port 12 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 40000 40733
string GDS_END 35677486
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 35412430
string LEFclass PAD
string LEFsymmetry X Y R90
<< end >>
