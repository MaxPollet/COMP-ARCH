magic
tech sky130A
magscale 1 2
timestamp 1681267127
<< nwell >>
rect -66 377 3138 897
<< pwell >>
rect 454 217 1974 283
rect 2623 217 3068 317
rect 4 43 3068 217
rect -26 -43 3098 43
<< locali >>
rect 112 235 178 430
rect 539 324 647 498
rect 613 126 647 324
rect 683 162 749 421
rect 1321 365 1692 399
rect 1658 259 1692 365
rect 1168 225 1692 259
rect 1168 126 1202 225
rect 613 92 1202 126
rect 1658 87 1692 225
rect 2291 253 2357 331
rect 2156 219 2357 253
rect 2156 87 2190 219
rect 1658 53 2190 87
rect 2980 133 3047 747
<< obsli1 >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 3007 831
rect 3041 797 3072 831
rect 126 735 244 741
rect 126 701 132 735
rect 166 701 204 735
rect 238 701 244 735
rect 22 505 88 691
rect 126 545 244 701
rect 280 727 568 761
rect 280 505 314 727
rect 22 471 314 505
rect 22 99 76 471
rect 248 371 314 471
rect 350 430 400 691
rect 448 568 498 691
rect 534 638 568 727
rect 604 735 670 741
rect 604 701 610 735
rect 644 701 670 735
rect 604 674 670 701
rect 706 727 1054 761
rect 706 638 740 727
rect 534 604 740 638
rect 776 568 810 691
rect 916 640 982 691
rect 448 534 810 568
rect 846 534 890 600
rect 776 498 810 534
rect 350 384 455 430
rect 350 199 404 384
rect 776 464 820 498
rect 112 113 302 199
rect 112 79 118 113
rect 152 79 190 113
rect 224 79 262 113
rect 296 79 302 113
rect 338 99 404 199
rect 440 113 558 249
rect 112 73 302 79
rect 440 79 446 113
rect 480 79 518 113
rect 552 79 558 113
rect 786 265 820 464
rect 856 430 890 534
rect 926 500 960 640
rect 1020 609 1054 727
rect 1090 735 1280 741
rect 1090 701 1096 735
rect 1130 701 1168 735
rect 1202 701 1240 735
rect 1274 701 1280 735
rect 1090 645 1280 701
rect 1316 727 1522 761
rect 1316 609 1350 727
rect 1020 600 1350 609
rect 996 575 1350 600
rect 996 536 1062 575
rect 1386 539 1452 691
rect 1488 655 1522 727
rect 1558 735 1748 751
rect 1558 701 1564 735
rect 1598 701 1636 735
rect 1670 701 1708 735
rect 1742 701 1748 735
rect 1558 691 1748 701
rect 1488 621 1850 655
rect 1098 505 1452 539
rect 1098 500 1132 505
rect 926 466 1132 500
rect 1714 469 1780 585
rect 856 384 1061 430
rect 995 285 1061 384
rect 1098 329 1132 466
rect 1168 435 1780 469
rect 1168 365 1234 435
rect 1098 295 1622 329
rect 786 165 840 265
rect 1098 249 1132 295
rect 930 215 1132 249
rect 930 165 996 215
rect 1432 113 1622 189
rect 440 73 558 79
rect 1432 79 1438 113
rect 1472 79 1510 113
rect 1544 79 1582 113
rect 1616 79 1622 113
rect 1432 73 1622 79
rect 1728 265 1780 435
rect 1816 351 1850 621
rect 1886 569 1936 751
rect 2097 735 2287 741
rect 2097 701 2103 735
rect 2137 701 2175 735
rect 2209 701 2247 735
rect 2281 701 2287 735
rect 1886 535 2061 569
rect 2097 535 2287 701
rect 2454 735 2633 741
rect 2488 701 2526 735
rect 2560 701 2598 735
rect 2632 701 2633 735
rect 2368 541 2418 635
rect 2454 577 2633 701
rect 2755 735 2944 747
rect 2755 701 2760 735
rect 2794 701 2832 735
rect 2866 701 2904 735
rect 2938 701 2944 735
rect 1925 387 1991 487
rect 2027 471 2061 535
rect 2368 507 2569 541
rect 2027 437 2499 471
rect 1816 317 2050 351
rect 1728 123 1794 265
rect 1886 157 1952 265
rect 1993 217 2050 317
rect 2086 157 2120 437
rect 2535 401 2569 507
rect 2161 367 2569 401
rect 2161 289 2227 367
rect 1886 123 2120 157
rect 2524 199 2569 367
rect 2669 401 2719 601
rect 2755 439 2944 701
rect 2669 335 2944 401
rect 2669 299 2711 335
rect 2645 199 2711 299
rect 2226 113 2416 183
rect 2226 79 2232 113
rect 2266 79 2304 113
rect 2338 79 2376 113
rect 2410 79 2416 113
rect 2524 99 2590 199
rect 2747 113 2937 299
rect 2226 73 2416 79
rect 2747 79 2753 113
rect 2787 79 2825 113
rect 2859 79 2897 113
rect 2931 79 2937 113
rect 2747 73 2937 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3072 17
<< obsli1c >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 2143 797 2177 831
rect 2239 797 2273 831
rect 2335 797 2369 831
rect 2431 797 2465 831
rect 2527 797 2561 831
rect 2623 797 2657 831
rect 2719 797 2753 831
rect 2815 797 2849 831
rect 2911 797 2945 831
rect 3007 797 3041 831
rect 132 701 166 735
rect 204 701 238 735
rect 610 701 644 735
rect 118 79 152 113
rect 190 79 224 113
rect 262 79 296 113
rect 446 79 480 113
rect 518 79 552 113
rect 1096 701 1130 735
rect 1168 701 1202 735
rect 1240 701 1274 735
rect 1564 701 1598 735
rect 1636 701 1670 735
rect 1708 701 1742 735
rect 1438 79 1472 113
rect 1510 79 1544 113
rect 1582 79 1616 113
rect 2103 701 2137 735
rect 2175 701 2209 735
rect 2247 701 2281 735
rect 2454 701 2488 735
rect 2526 701 2560 735
rect 2598 701 2632 735
rect 2760 701 2794 735
rect 2832 701 2866 735
rect 2904 701 2938 735
rect 2232 79 2266 113
rect 2304 79 2338 113
rect 2376 79 2410 113
rect 2753 79 2787 113
rect 2825 79 2859 113
rect 2897 79 2931 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
<< metal1 >>
rect 0 831 3072 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 3007 831
rect 3041 797 3072 831
rect 0 791 3072 797
rect 0 735 3072 763
rect 0 701 132 735
rect 166 701 204 735
rect 238 701 610 735
rect 644 701 1096 735
rect 1130 701 1168 735
rect 1202 701 1240 735
rect 1274 701 1564 735
rect 1598 701 1636 735
rect 1670 701 1708 735
rect 1742 701 2103 735
rect 2137 701 2175 735
rect 2209 701 2247 735
rect 2281 701 2454 735
rect 2488 701 2526 735
rect 2560 701 2598 735
rect 2632 701 2760 735
rect 2794 701 2832 735
rect 2866 701 2904 735
rect 2938 701 3072 735
rect 0 689 3072 701
rect 0 113 3072 125
rect 0 79 118 113
rect 152 79 190 113
rect 224 79 262 113
rect 296 79 446 113
rect 480 79 518 113
rect 552 79 1438 113
rect 1472 79 1510 113
rect 1544 79 1582 113
rect 1616 79 2232 113
rect 2266 79 2304 113
rect 2338 79 2376 113
rect 2410 79 2753 113
rect 2787 79 2825 113
rect 2859 79 2897 113
rect 2931 79 3072 113
rect 0 51 3072 79
rect 0 17 3072 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3072 17
rect 0 -23 3072 -17
<< obsm1 >>
rect 403 421 461 430
rect 883 421 941 430
rect 1939 421 1997 430
rect 403 393 1997 421
rect 403 384 461 393
rect 883 384 941 393
rect 1939 384 1997 393
<< labels >>
rlabel locali s 112 235 178 430 6 CLK
port 1 nsew clock input
rlabel locali s 683 162 749 421 6 D
port 2 nsew signal input
rlabel locali s 1658 53 2190 87 6 RESET_B
port 3 nsew signal input
rlabel locali s 2156 87 2190 219 6 RESET_B
port 3 nsew signal input
rlabel locali s 2156 219 2357 253 6 RESET_B
port 3 nsew signal input
rlabel locali s 1658 87 1692 225 6 RESET_B
port 3 nsew signal input
rlabel locali s 613 92 1202 126 6 RESET_B
port 3 nsew signal input
rlabel locali s 1168 126 1202 225 6 RESET_B
port 3 nsew signal input
rlabel locali s 2291 253 2357 331 6 RESET_B
port 3 nsew signal input
rlabel locali s 1168 225 1692 259 6 RESET_B
port 3 nsew signal input
rlabel locali s 1658 259 1692 365 6 RESET_B
port 3 nsew signal input
rlabel locali s 613 126 647 324 6 RESET_B
port 3 nsew signal input
rlabel locali s 1321 365 1692 399 6 RESET_B
port 3 nsew signal input
rlabel locali s 539 324 647 498 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 0 51 3072 125 6 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 -23 3072 23 8 VNB
port 5 nsew ground bidirectional
rlabel pwell s -26 -43 3098 43 8 VNB
port 5 nsew ground bidirectional
rlabel pwell s 4 43 3068 217 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 2623 217 3068 317 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 454 217 1974 283 6 VNB
port 5 nsew ground bidirectional
rlabel metal1 s 0 791 3072 837 6 VPB
port 6 nsew power bidirectional
rlabel nwell s -66 377 3138 897 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 689 3072 763 6 VPWR
port 7 nsew power bidirectional
rlabel locali s 2980 133 3047 747 6 Q
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 3072 814
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 948166
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 919000
<< end >>
