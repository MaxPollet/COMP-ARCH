magic
tech sky130A
magscale 1 2
timestamp 1681267127
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 1 21 813 203
rect 29 -17 63 21
<< locali >>
rect 17 291 122 493
rect 17 177 71 291
rect 255 215 339 257
rect 373 215 439 478
rect 481 215 547 478
rect 581 215 655 478
rect 697 215 799 265
rect 17 51 85 177
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 169 383 235 527
rect 269 349 319 493
rect 169 291 319 349
rect 169 257 221 291
rect 105 215 221 257
rect 721 303 787 527
rect 147 181 221 215
rect 147 143 297 181
rect 143 17 177 109
rect 231 54 297 143
rect 331 147 791 181
rect 331 83 365 147
rect 410 17 476 109
rect 516 51 582 147
rect 625 17 691 109
rect 725 51 791 147
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
rlabel locali s 697 215 799 265 6 A1
port 1 nsew signal input
rlabel locali s 581 215 655 478 6 A2
port 2 nsew signal input
rlabel locali s 481 215 547 478 6 A3
port 3 nsew signal input
rlabel locali s 373 215 439 478 6 A4
port 4 nsew signal input
rlabel locali s 255 215 339 257 6 B1
port 5 nsew signal input
rlabel metal1 s 0 -48 828 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 1 21 813 203 6 VNB
port 7 nsew ground bidirectional
rlabel nwell s -38 261 866 582 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 496 828 592 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 17 51 85 177 6 X
port 10 nsew signal output
rlabel locali s 17 177 71 291 6 X
port 10 nsew signal output
rlabel locali s 17 291 122 493 6 X
port 10 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 828 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1521832
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1513678
<< end >>
