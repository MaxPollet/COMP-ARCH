magic
tech sky130A
magscale 1 2
timestamp 1681267127
<< pwell >>
rect 10 66 1014 1128
<< mvnmos >>
rect 228 92 328 1102
rect 384 92 484 1102
rect 540 92 640 1102
rect 696 92 796 1102
<< mvndiff >>
rect 172 1090 228 1102
rect 172 1056 183 1090
rect 217 1056 228 1090
rect 172 1022 228 1056
rect 172 988 183 1022
rect 217 988 228 1022
rect 172 954 228 988
rect 172 920 183 954
rect 217 920 228 954
rect 172 886 228 920
rect 172 852 183 886
rect 217 852 228 886
rect 172 818 228 852
rect 172 784 183 818
rect 217 784 228 818
rect 172 750 228 784
rect 172 716 183 750
rect 217 716 228 750
rect 172 682 228 716
rect 172 648 183 682
rect 217 648 228 682
rect 172 614 228 648
rect 172 580 183 614
rect 217 580 228 614
rect 172 546 228 580
rect 172 512 183 546
rect 217 512 228 546
rect 172 478 228 512
rect 172 444 183 478
rect 217 444 228 478
rect 172 410 228 444
rect 172 376 183 410
rect 217 376 228 410
rect 172 342 228 376
rect 172 308 183 342
rect 217 308 228 342
rect 172 274 228 308
rect 172 240 183 274
rect 217 240 228 274
rect 172 206 228 240
rect 172 172 183 206
rect 217 172 228 206
rect 172 138 228 172
rect 172 104 183 138
rect 217 104 228 138
rect 172 92 228 104
rect 328 1090 384 1102
rect 328 1056 339 1090
rect 373 1056 384 1090
rect 328 1022 384 1056
rect 328 988 339 1022
rect 373 988 384 1022
rect 328 954 384 988
rect 328 920 339 954
rect 373 920 384 954
rect 328 886 384 920
rect 328 852 339 886
rect 373 852 384 886
rect 328 818 384 852
rect 328 784 339 818
rect 373 784 384 818
rect 328 750 384 784
rect 328 716 339 750
rect 373 716 384 750
rect 328 682 384 716
rect 328 648 339 682
rect 373 648 384 682
rect 328 614 384 648
rect 328 580 339 614
rect 373 580 384 614
rect 328 546 384 580
rect 328 512 339 546
rect 373 512 384 546
rect 328 478 384 512
rect 328 444 339 478
rect 373 444 384 478
rect 328 410 384 444
rect 328 376 339 410
rect 373 376 384 410
rect 328 342 384 376
rect 328 308 339 342
rect 373 308 384 342
rect 328 274 384 308
rect 328 240 339 274
rect 373 240 384 274
rect 328 206 384 240
rect 328 172 339 206
rect 373 172 384 206
rect 328 138 384 172
rect 328 104 339 138
rect 373 104 384 138
rect 328 92 384 104
rect 484 1090 540 1102
rect 484 1056 495 1090
rect 529 1056 540 1090
rect 484 1022 540 1056
rect 484 988 495 1022
rect 529 988 540 1022
rect 484 954 540 988
rect 484 920 495 954
rect 529 920 540 954
rect 484 886 540 920
rect 484 852 495 886
rect 529 852 540 886
rect 484 818 540 852
rect 484 784 495 818
rect 529 784 540 818
rect 484 750 540 784
rect 484 716 495 750
rect 529 716 540 750
rect 484 682 540 716
rect 484 648 495 682
rect 529 648 540 682
rect 484 614 540 648
rect 484 580 495 614
rect 529 580 540 614
rect 484 546 540 580
rect 484 512 495 546
rect 529 512 540 546
rect 484 478 540 512
rect 484 444 495 478
rect 529 444 540 478
rect 484 410 540 444
rect 484 376 495 410
rect 529 376 540 410
rect 484 342 540 376
rect 484 308 495 342
rect 529 308 540 342
rect 484 274 540 308
rect 484 240 495 274
rect 529 240 540 274
rect 484 206 540 240
rect 484 172 495 206
rect 529 172 540 206
rect 484 138 540 172
rect 484 104 495 138
rect 529 104 540 138
rect 484 92 540 104
rect 640 1090 696 1102
rect 640 1056 651 1090
rect 685 1056 696 1090
rect 640 1022 696 1056
rect 640 988 651 1022
rect 685 988 696 1022
rect 640 954 696 988
rect 640 920 651 954
rect 685 920 696 954
rect 640 886 696 920
rect 640 852 651 886
rect 685 852 696 886
rect 640 818 696 852
rect 640 784 651 818
rect 685 784 696 818
rect 640 750 696 784
rect 640 716 651 750
rect 685 716 696 750
rect 640 682 696 716
rect 640 648 651 682
rect 685 648 696 682
rect 640 614 696 648
rect 640 580 651 614
rect 685 580 696 614
rect 640 546 696 580
rect 640 512 651 546
rect 685 512 696 546
rect 640 478 696 512
rect 640 444 651 478
rect 685 444 696 478
rect 640 410 696 444
rect 640 376 651 410
rect 685 376 696 410
rect 640 342 696 376
rect 640 308 651 342
rect 685 308 696 342
rect 640 274 696 308
rect 640 240 651 274
rect 685 240 696 274
rect 640 206 696 240
rect 640 172 651 206
rect 685 172 696 206
rect 640 138 696 172
rect 640 104 651 138
rect 685 104 696 138
rect 640 92 696 104
rect 796 1090 852 1102
rect 796 1056 807 1090
rect 841 1056 852 1090
rect 796 1022 852 1056
rect 796 988 807 1022
rect 841 988 852 1022
rect 796 954 852 988
rect 796 920 807 954
rect 841 920 852 954
rect 796 886 852 920
rect 796 852 807 886
rect 841 852 852 886
rect 796 818 852 852
rect 796 784 807 818
rect 841 784 852 818
rect 796 750 852 784
rect 796 716 807 750
rect 841 716 852 750
rect 796 682 852 716
rect 796 648 807 682
rect 841 648 852 682
rect 796 614 852 648
rect 796 580 807 614
rect 841 580 852 614
rect 796 546 852 580
rect 796 512 807 546
rect 841 512 852 546
rect 796 478 852 512
rect 796 444 807 478
rect 841 444 852 478
rect 796 410 852 444
rect 796 376 807 410
rect 841 376 852 410
rect 796 342 852 376
rect 796 308 807 342
rect 841 308 852 342
rect 796 274 852 308
rect 796 240 807 274
rect 841 240 852 274
rect 796 206 852 240
rect 796 172 807 206
rect 841 172 852 206
rect 796 138 852 172
rect 796 104 807 138
rect 841 104 852 138
rect 796 92 852 104
<< mvndiffc >>
rect 183 1056 217 1090
rect 183 988 217 1022
rect 183 920 217 954
rect 183 852 217 886
rect 183 784 217 818
rect 183 716 217 750
rect 183 648 217 682
rect 183 580 217 614
rect 183 512 217 546
rect 183 444 217 478
rect 183 376 217 410
rect 183 308 217 342
rect 183 240 217 274
rect 183 172 217 206
rect 183 104 217 138
rect 339 1056 373 1090
rect 339 988 373 1022
rect 339 920 373 954
rect 339 852 373 886
rect 339 784 373 818
rect 339 716 373 750
rect 339 648 373 682
rect 339 580 373 614
rect 339 512 373 546
rect 339 444 373 478
rect 339 376 373 410
rect 339 308 373 342
rect 339 240 373 274
rect 339 172 373 206
rect 339 104 373 138
rect 495 1056 529 1090
rect 495 988 529 1022
rect 495 920 529 954
rect 495 852 529 886
rect 495 784 529 818
rect 495 716 529 750
rect 495 648 529 682
rect 495 580 529 614
rect 495 512 529 546
rect 495 444 529 478
rect 495 376 529 410
rect 495 308 529 342
rect 495 240 529 274
rect 495 172 529 206
rect 495 104 529 138
rect 651 1056 685 1090
rect 651 988 685 1022
rect 651 920 685 954
rect 651 852 685 886
rect 651 784 685 818
rect 651 716 685 750
rect 651 648 685 682
rect 651 580 685 614
rect 651 512 685 546
rect 651 444 685 478
rect 651 376 685 410
rect 651 308 685 342
rect 651 240 685 274
rect 651 172 685 206
rect 651 104 685 138
rect 807 1056 841 1090
rect 807 988 841 1022
rect 807 920 841 954
rect 807 852 841 886
rect 807 784 841 818
rect 807 716 841 750
rect 807 648 841 682
rect 807 580 841 614
rect 807 512 841 546
rect 807 444 841 478
rect 807 376 841 410
rect 807 308 841 342
rect 807 240 841 274
rect 807 172 841 206
rect 807 104 841 138
<< mvpsubdiff >>
rect 36 1056 94 1102
rect 36 1022 48 1056
rect 82 1022 94 1056
rect 36 988 94 1022
rect 36 954 48 988
rect 82 954 94 988
rect 36 920 94 954
rect 36 886 48 920
rect 82 886 94 920
rect 36 852 94 886
rect 36 818 48 852
rect 82 818 94 852
rect 36 784 94 818
rect 36 750 48 784
rect 82 750 94 784
rect 36 716 94 750
rect 36 682 48 716
rect 82 682 94 716
rect 36 648 94 682
rect 36 614 48 648
rect 82 614 94 648
rect 36 580 94 614
rect 36 546 48 580
rect 82 546 94 580
rect 36 512 94 546
rect 36 478 48 512
rect 82 478 94 512
rect 36 444 94 478
rect 36 410 48 444
rect 82 410 94 444
rect 36 376 94 410
rect 36 342 48 376
rect 82 342 94 376
rect 36 308 94 342
rect 36 274 48 308
rect 82 274 94 308
rect 36 240 94 274
rect 36 206 48 240
rect 82 206 94 240
rect 36 172 94 206
rect 36 138 48 172
rect 82 138 94 172
rect 36 92 94 138
rect 930 1056 988 1102
rect 930 1022 942 1056
rect 976 1022 988 1056
rect 930 988 988 1022
rect 930 954 942 988
rect 976 954 988 988
rect 930 920 988 954
rect 930 886 942 920
rect 976 886 988 920
rect 930 852 988 886
rect 930 818 942 852
rect 976 818 988 852
rect 930 784 988 818
rect 930 750 942 784
rect 976 750 988 784
rect 930 716 988 750
rect 930 682 942 716
rect 976 682 988 716
rect 930 648 988 682
rect 930 614 942 648
rect 976 614 988 648
rect 930 580 988 614
rect 930 546 942 580
rect 976 546 988 580
rect 930 512 988 546
rect 930 478 942 512
rect 976 478 988 512
rect 930 444 988 478
rect 930 410 942 444
rect 976 410 988 444
rect 930 376 988 410
rect 930 342 942 376
rect 976 342 988 376
rect 930 308 988 342
rect 930 274 942 308
rect 976 274 988 308
rect 930 240 988 274
rect 930 206 942 240
rect 976 206 988 240
rect 930 172 988 206
rect 930 138 942 172
rect 976 138 988 172
rect 930 92 988 138
<< mvpsubdiffcont >>
rect 48 1022 82 1056
rect 48 954 82 988
rect 48 886 82 920
rect 48 818 82 852
rect 48 750 82 784
rect 48 682 82 716
rect 48 614 82 648
rect 48 546 82 580
rect 48 478 82 512
rect 48 410 82 444
rect 48 342 82 376
rect 48 274 82 308
rect 48 206 82 240
rect 48 138 82 172
rect 942 1022 976 1056
rect 942 954 976 988
rect 942 886 976 920
rect 942 818 976 852
rect 942 750 976 784
rect 942 682 976 716
rect 942 614 976 648
rect 942 546 976 580
rect 942 478 976 512
rect 942 410 976 444
rect 942 342 976 376
rect 942 274 976 308
rect 942 206 976 240
rect 942 138 976 172
<< poly >>
rect 207 1174 817 1194
rect 207 1140 223 1174
rect 257 1140 291 1174
rect 325 1140 359 1174
rect 393 1140 427 1174
rect 461 1140 495 1174
rect 529 1140 563 1174
rect 597 1140 631 1174
rect 665 1140 699 1174
rect 733 1140 767 1174
rect 801 1140 817 1174
rect 207 1124 817 1140
rect 228 1102 328 1124
rect 384 1102 484 1124
rect 540 1102 640 1124
rect 696 1102 796 1124
rect 228 70 328 92
rect 384 70 484 92
rect 540 70 640 92
rect 696 70 796 92
rect 207 54 817 70
rect 207 20 223 54
rect 257 20 291 54
rect 325 20 359 54
rect 393 20 427 54
rect 461 20 495 54
rect 529 20 563 54
rect 597 20 631 54
rect 665 20 699 54
rect 733 20 767 54
rect 801 20 817 54
rect 207 0 817 20
<< polycont >>
rect 223 1140 257 1174
rect 291 1140 325 1174
rect 359 1140 393 1174
rect 427 1140 461 1174
rect 495 1140 529 1174
rect 563 1140 597 1174
rect 631 1140 665 1174
rect 699 1140 733 1174
rect 767 1140 801 1174
rect 223 20 257 54
rect 291 20 325 54
rect 359 20 393 54
rect 427 20 461 54
rect 495 20 529 54
rect 563 20 597 54
rect 631 20 665 54
rect 699 20 733 54
rect 767 20 801 54
<< locali >>
rect 207 1140 223 1174
rect 277 1140 291 1174
rect 349 1140 359 1174
rect 421 1140 427 1174
rect 493 1140 495 1174
rect 529 1140 531 1174
rect 597 1140 603 1174
rect 665 1140 675 1174
rect 733 1140 747 1174
rect 801 1140 817 1174
rect 183 1090 217 1106
rect 48 1010 82 1022
rect 48 938 82 954
rect 48 866 82 886
rect 48 794 82 818
rect 48 722 82 750
rect 48 650 82 682
rect 48 580 82 614
rect 48 512 82 544
rect 48 444 82 472
rect 48 376 82 400
rect 48 308 82 328
rect 48 240 82 256
rect 48 172 82 184
rect 183 1022 217 1048
rect 183 954 217 976
rect 183 886 217 904
rect 183 818 217 832
rect 183 750 217 760
rect 183 682 217 688
rect 183 614 217 616
rect 183 578 217 580
rect 183 506 217 512
rect 183 434 217 444
rect 183 362 217 376
rect 183 290 217 308
rect 183 218 217 240
rect 183 146 217 172
rect 183 88 217 104
rect 339 1090 373 1106
rect 339 1022 373 1048
rect 339 954 373 976
rect 339 886 373 904
rect 339 818 373 832
rect 339 750 373 760
rect 339 682 373 688
rect 339 614 373 616
rect 339 578 373 580
rect 339 506 373 512
rect 339 434 373 444
rect 339 362 373 376
rect 339 290 373 308
rect 339 218 373 240
rect 339 146 373 172
rect 339 88 373 104
rect 495 1090 529 1106
rect 495 1022 529 1048
rect 495 954 529 976
rect 495 886 529 904
rect 495 818 529 832
rect 495 750 529 760
rect 495 682 529 688
rect 495 614 529 616
rect 495 578 529 580
rect 495 506 529 512
rect 495 434 529 444
rect 495 362 529 376
rect 495 290 529 308
rect 495 218 529 240
rect 495 146 529 172
rect 495 88 529 104
rect 651 1090 685 1106
rect 651 1022 685 1048
rect 651 954 685 976
rect 651 886 685 904
rect 651 818 685 832
rect 651 750 685 760
rect 651 682 685 688
rect 651 614 685 616
rect 651 578 685 580
rect 651 506 685 512
rect 651 434 685 444
rect 651 362 685 376
rect 651 290 685 308
rect 651 218 685 240
rect 651 146 685 172
rect 651 88 685 104
rect 807 1090 841 1106
rect 807 1022 841 1048
rect 807 954 841 976
rect 807 886 841 904
rect 807 818 841 832
rect 807 750 841 760
rect 807 682 841 688
rect 807 614 841 616
rect 807 578 841 580
rect 807 506 841 512
rect 807 434 841 444
rect 807 362 841 376
rect 807 290 841 308
rect 807 218 841 240
rect 807 146 841 172
rect 942 1010 976 1022
rect 942 938 976 954
rect 942 866 976 886
rect 942 794 976 818
rect 942 722 976 750
rect 942 650 976 682
rect 942 580 976 614
rect 942 512 976 544
rect 942 444 976 472
rect 942 376 976 400
rect 942 308 976 328
rect 942 240 976 256
rect 942 172 976 184
rect 807 88 841 104
rect 207 20 223 54
rect 277 20 291 54
rect 349 20 359 54
rect 421 20 427 54
rect 493 20 495 54
rect 529 20 531 54
rect 597 20 603 54
rect 665 20 675 54
rect 733 20 747 54
rect 801 20 817 54
<< viali >>
rect 243 1140 257 1174
rect 257 1140 277 1174
rect 315 1140 325 1174
rect 325 1140 349 1174
rect 387 1140 393 1174
rect 393 1140 421 1174
rect 459 1140 461 1174
rect 461 1140 493 1174
rect 531 1140 563 1174
rect 563 1140 565 1174
rect 603 1140 631 1174
rect 631 1140 637 1174
rect 675 1140 699 1174
rect 699 1140 709 1174
rect 747 1140 767 1174
rect 767 1140 781 1174
rect 48 1056 82 1082
rect 48 1048 82 1056
rect 48 988 82 1010
rect 48 976 82 988
rect 48 920 82 938
rect 48 904 82 920
rect 48 852 82 866
rect 48 832 82 852
rect 48 784 82 794
rect 48 760 82 784
rect 48 716 82 722
rect 48 688 82 716
rect 48 648 82 650
rect 48 616 82 648
rect 48 546 82 578
rect 48 544 82 546
rect 48 478 82 506
rect 48 472 82 478
rect 48 410 82 434
rect 48 400 82 410
rect 48 342 82 362
rect 48 328 82 342
rect 48 274 82 290
rect 48 256 82 274
rect 48 206 82 218
rect 48 184 82 206
rect 48 138 82 146
rect 48 112 82 138
rect 183 1056 217 1082
rect 183 1048 217 1056
rect 183 988 217 1010
rect 183 976 217 988
rect 183 920 217 938
rect 183 904 217 920
rect 183 852 217 866
rect 183 832 217 852
rect 183 784 217 794
rect 183 760 217 784
rect 183 716 217 722
rect 183 688 217 716
rect 183 648 217 650
rect 183 616 217 648
rect 183 546 217 578
rect 183 544 217 546
rect 183 478 217 506
rect 183 472 217 478
rect 183 410 217 434
rect 183 400 217 410
rect 183 342 217 362
rect 183 328 217 342
rect 183 274 217 290
rect 183 256 217 274
rect 183 206 217 218
rect 183 184 217 206
rect 183 138 217 146
rect 183 112 217 138
rect 339 1056 373 1082
rect 339 1048 373 1056
rect 339 988 373 1010
rect 339 976 373 988
rect 339 920 373 938
rect 339 904 373 920
rect 339 852 373 866
rect 339 832 373 852
rect 339 784 373 794
rect 339 760 373 784
rect 339 716 373 722
rect 339 688 373 716
rect 339 648 373 650
rect 339 616 373 648
rect 339 546 373 578
rect 339 544 373 546
rect 339 478 373 506
rect 339 472 373 478
rect 339 410 373 434
rect 339 400 373 410
rect 339 342 373 362
rect 339 328 373 342
rect 339 274 373 290
rect 339 256 373 274
rect 339 206 373 218
rect 339 184 373 206
rect 339 138 373 146
rect 339 112 373 138
rect 495 1056 529 1082
rect 495 1048 529 1056
rect 495 988 529 1010
rect 495 976 529 988
rect 495 920 529 938
rect 495 904 529 920
rect 495 852 529 866
rect 495 832 529 852
rect 495 784 529 794
rect 495 760 529 784
rect 495 716 529 722
rect 495 688 529 716
rect 495 648 529 650
rect 495 616 529 648
rect 495 546 529 578
rect 495 544 529 546
rect 495 478 529 506
rect 495 472 529 478
rect 495 410 529 434
rect 495 400 529 410
rect 495 342 529 362
rect 495 328 529 342
rect 495 274 529 290
rect 495 256 529 274
rect 495 206 529 218
rect 495 184 529 206
rect 495 138 529 146
rect 495 112 529 138
rect 651 1056 685 1082
rect 651 1048 685 1056
rect 651 988 685 1010
rect 651 976 685 988
rect 651 920 685 938
rect 651 904 685 920
rect 651 852 685 866
rect 651 832 685 852
rect 651 784 685 794
rect 651 760 685 784
rect 651 716 685 722
rect 651 688 685 716
rect 651 648 685 650
rect 651 616 685 648
rect 651 546 685 578
rect 651 544 685 546
rect 651 478 685 506
rect 651 472 685 478
rect 651 410 685 434
rect 651 400 685 410
rect 651 342 685 362
rect 651 328 685 342
rect 651 274 685 290
rect 651 256 685 274
rect 651 206 685 218
rect 651 184 685 206
rect 651 138 685 146
rect 651 112 685 138
rect 807 1056 841 1082
rect 807 1048 841 1056
rect 807 988 841 1010
rect 807 976 841 988
rect 807 920 841 938
rect 807 904 841 920
rect 807 852 841 866
rect 807 832 841 852
rect 807 784 841 794
rect 807 760 841 784
rect 807 716 841 722
rect 807 688 841 716
rect 807 648 841 650
rect 807 616 841 648
rect 807 546 841 578
rect 807 544 841 546
rect 807 478 841 506
rect 807 472 841 478
rect 807 410 841 434
rect 807 400 841 410
rect 807 342 841 362
rect 807 328 841 342
rect 807 274 841 290
rect 807 256 841 274
rect 807 206 841 218
rect 807 184 841 206
rect 807 138 841 146
rect 807 112 841 138
rect 942 1056 976 1082
rect 942 1048 976 1056
rect 942 988 976 1010
rect 942 976 976 988
rect 942 920 976 938
rect 942 904 976 920
rect 942 852 976 866
rect 942 832 976 852
rect 942 784 976 794
rect 942 760 976 784
rect 942 716 976 722
rect 942 688 976 716
rect 942 648 976 650
rect 942 616 976 648
rect 942 546 976 578
rect 942 544 976 546
rect 942 478 976 506
rect 942 472 976 478
rect 942 410 976 434
rect 942 400 976 410
rect 942 342 976 362
rect 942 328 976 342
rect 942 274 976 290
rect 942 256 976 274
rect 942 206 976 218
rect 942 184 976 206
rect 942 138 976 146
rect 942 112 976 138
rect 243 20 257 54
rect 257 20 277 54
rect 315 20 325 54
rect 325 20 349 54
rect 387 20 393 54
rect 393 20 421 54
rect 459 20 461 54
rect 461 20 493 54
rect 531 20 563 54
rect 563 20 565 54
rect 603 20 631 54
rect 631 20 637 54
rect 675 20 699 54
rect 699 20 709 54
rect 747 20 767 54
rect 767 20 781 54
<< metal1 >>
rect 231 1174 793 1194
rect 231 1140 243 1174
rect 277 1140 315 1174
rect 349 1140 387 1174
rect 421 1140 459 1174
rect 493 1140 531 1174
rect 565 1140 603 1174
rect 637 1140 675 1174
rect 709 1140 747 1174
rect 781 1140 793 1174
rect 231 1128 793 1140
rect 36 1082 95 1094
rect 36 1048 48 1082
rect 82 1048 95 1082
rect 36 1010 95 1048
rect 36 976 48 1010
rect 82 976 95 1010
rect 36 938 95 976
rect 36 904 48 938
rect 82 904 95 938
rect 36 866 95 904
rect 36 832 48 866
rect 82 832 95 866
rect 36 794 95 832
rect 36 760 48 794
rect 82 760 95 794
rect 36 722 95 760
rect 36 688 48 722
rect 82 688 95 722
rect 36 650 95 688
rect 36 616 48 650
rect 82 616 95 650
rect 36 578 95 616
rect 36 544 48 578
rect 82 544 95 578
rect 36 506 95 544
rect 36 472 48 506
rect 82 472 95 506
rect 36 434 95 472
rect 36 400 48 434
rect 82 400 95 434
rect 36 362 95 400
rect 36 328 48 362
rect 82 328 95 362
rect 36 290 95 328
rect 36 256 48 290
rect 82 256 95 290
rect 36 218 95 256
rect 36 184 48 218
rect 82 184 95 218
rect 36 146 95 184
rect 36 112 48 146
rect 82 112 95 146
rect 36 100 95 112
rect 174 1082 226 1094
rect 174 1048 183 1082
rect 217 1048 226 1082
rect 174 1010 226 1048
rect 174 976 183 1010
rect 217 976 226 1010
rect 174 938 226 976
rect 174 904 183 938
rect 217 904 226 938
rect 174 866 226 904
rect 174 832 183 866
rect 217 832 226 866
rect 174 794 226 832
rect 174 760 183 794
rect 217 760 226 794
rect 174 722 226 760
rect 174 688 183 722
rect 217 688 226 722
rect 174 650 226 688
rect 174 616 183 650
rect 217 616 226 650
rect 174 578 226 616
rect 174 544 183 578
rect 217 544 226 578
rect 174 542 226 544
rect 174 478 183 490
rect 217 478 226 490
rect 174 414 183 426
rect 217 414 226 426
rect 174 350 183 362
rect 217 350 226 362
rect 174 290 226 298
rect 174 286 183 290
rect 217 286 226 290
rect 174 222 226 234
rect 174 158 226 170
rect 174 100 226 106
rect 330 1088 382 1094
rect 330 1024 382 1036
rect 330 960 382 972
rect 330 904 339 908
rect 373 904 382 908
rect 330 896 382 904
rect 330 832 339 844
rect 373 832 382 844
rect 330 768 339 780
rect 373 768 382 780
rect 330 704 339 716
rect 373 704 382 716
rect 330 650 382 652
rect 330 616 339 650
rect 373 616 382 650
rect 330 578 382 616
rect 330 544 339 578
rect 373 544 382 578
rect 330 506 382 544
rect 330 472 339 506
rect 373 472 382 506
rect 330 434 382 472
rect 330 400 339 434
rect 373 400 382 434
rect 330 362 382 400
rect 330 328 339 362
rect 373 328 382 362
rect 330 290 382 328
rect 330 256 339 290
rect 373 256 382 290
rect 330 218 382 256
rect 330 184 339 218
rect 373 184 382 218
rect 330 146 382 184
rect 330 112 339 146
rect 373 112 382 146
rect 330 100 382 112
rect 486 1082 538 1094
rect 486 1048 495 1082
rect 529 1048 538 1082
rect 486 1010 538 1048
rect 486 976 495 1010
rect 529 976 538 1010
rect 486 938 538 976
rect 486 904 495 938
rect 529 904 538 938
rect 486 866 538 904
rect 486 832 495 866
rect 529 832 538 866
rect 486 794 538 832
rect 486 760 495 794
rect 529 760 538 794
rect 486 722 538 760
rect 486 688 495 722
rect 529 688 538 722
rect 486 650 538 688
rect 486 616 495 650
rect 529 616 538 650
rect 486 578 538 616
rect 486 544 495 578
rect 529 544 538 578
rect 486 542 538 544
rect 486 478 495 490
rect 529 478 538 490
rect 486 414 495 426
rect 529 414 538 426
rect 486 350 495 362
rect 529 350 538 362
rect 486 290 538 298
rect 486 286 495 290
rect 529 286 538 290
rect 486 222 538 234
rect 486 158 538 170
rect 486 100 538 106
rect 642 1088 694 1094
rect 642 1024 694 1036
rect 642 960 694 972
rect 642 904 651 908
rect 685 904 694 908
rect 642 896 694 904
rect 642 832 651 844
rect 685 832 694 844
rect 642 768 651 780
rect 685 768 694 780
rect 642 704 651 716
rect 685 704 694 716
rect 642 650 694 652
rect 642 616 651 650
rect 685 616 694 650
rect 642 578 694 616
rect 642 544 651 578
rect 685 544 694 578
rect 642 506 694 544
rect 642 472 651 506
rect 685 472 694 506
rect 642 434 694 472
rect 642 400 651 434
rect 685 400 694 434
rect 642 362 694 400
rect 642 328 651 362
rect 685 328 694 362
rect 642 290 694 328
rect 642 256 651 290
rect 685 256 694 290
rect 642 218 694 256
rect 642 184 651 218
rect 685 184 694 218
rect 642 146 694 184
rect 642 112 651 146
rect 685 112 694 146
rect 642 100 694 112
rect 798 1082 850 1094
rect 798 1048 807 1082
rect 841 1048 850 1082
rect 798 1010 850 1048
rect 798 976 807 1010
rect 841 976 850 1010
rect 798 938 850 976
rect 798 904 807 938
rect 841 904 850 938
rect 798 866 850 904
rect 798 832 807 866
rect 841 832 850 866
rect 798 794 850 832
rect 798 760 807 794
rect 841 760 850 794
rect 798 722 850 760
rect 798 688 807 722
rect 841 688 850 722
rect 798 650 850 688
rect 798 616 807 650
rect 841 616 850 650
rect 798 578 850 616
rect 798 544 807 578
rect 841 544 850 578
rect 798 542 850 544
rect 798 478 807 490
rect 841 478 850 490
rect 798 414 807 426
rect 841 414 850 426
rect 798 350 807 362
rect 841 350 850 362
rect 798 290 850 298
rect 798 286 807 290
rect 841 286 850 290
rect 798 222 850 234
rect 798 158 850 170
rect 798 100 850 106
rect 930 1082 989 1094
rect 930 1048 942 1082
rect 976 1048 989 1082
rect 930 1010 989 1048
rect 930 976 942 1010
rect 976 976 989 1010
rect 930 938 989 976
rect 930 904 942 938
rect 976 904 989 938
rect 930 866 989 904
rect 930 832 942 866
rect 976 832 989 866
rect 930 794 989 832
rect 930 760 942 794
rect 976 760 989 794
rect 930 722 989 760
rect 930 688 942 722
rect 976 688 989 722
rect 930 650 989 688
rect 930 616 942 650
rect 976 616 989 650
rect 930 578 989 616
rect 930 544 942 578
rect 976 544 989 578
rect 930 506 989 544
rect 930 472 942 506
rect 976 472 989 506
rect 930 434 989 472
rect 930 400 942 434
rect 976 400 989 434
rect 930 362 989 400
rect 930 328 942 362
rect 976 328 989 362
rect 930 290 989 328
rect 930 256 942 290
rect 976 256 989 290
rect 930 218 989 256
rect 930 184 942 218
rect 976 184 989 218
rect 930 146 989 184
rect 930 112 942 146
rect 976 112 989 146
rect 930 100 989 112
rect 231 54 793 66
rect 231 20 243 54
rect 277 20 315 54
rect 349 20 387 54
rect 421 20 459 54
rect 493 20 531 54
rect 565 20 603 54
rect 637 20 675 54
rect 709 20 747 54
rect 781 20 793 54
rect 231 0 793 20
<< via1 >>
rect 174 506 226 542
rect 174 490 183 506
rect 183 490 217 506
rect 217 490 226 506
rect 174 472 183 478
rect 183 472 217 478
rect 217 472 226 478
rect 174 434 226 472
rect 174 426 183 434
rect 183 426 217 434
rect 217 426 226 434
rect 174 400 183 414
rect 183 400 217 414
rect 217 400 226 414
rect 174 362 226 400
rect 174 328 183 350
rect 183 328 217 350
rect 217 328 226 350
rect 174 298 226 328
rect 174 256 183 286
rect 183 256 217 286
rect 217 256 226 286
rect 174 234 226 256
rect 174 218 226 222
rect 174 184 183 218
rect 183 184 217 218
rect 217 184 226 218
rect 174 170 226 184
rect 174 146 226 158
rect 174 112 183 146
rect 183 112 217 146
rect 217 112 226 146
rect 174 106 226 112
rect 330 1082 382 1088
rect 330 1048 339 1082
rect 339 1048 373 1082
rect 373 1048 382 1082
rect 330 1036 382 1048
rect 330 1010 382 1024
rect 330 976 339 1010
rect 339 976 373 1010
rect 373 976 382 1010
rect 330 972 382 976
rect 330 938 382 960
rect 330 908 339 938
rect 339 908 373 938
rect 373 908 382 938
rect 330 866 382 896
rect 330 844 339 866
rect 339 844 373 866
rect 373 844 382 866
rect 330 794 382 832
rect 330 780 339 794
rect 339 780 373 794
rect 373 780 382 794
rect 330 760 339 768
rect 339 760 373 768
rect 373 760 382 768
rect 330 722 382 760
rect 330 716 339 722
rect 339 716 373 722
rect 373 716 382 722
rect 330 688 339 704
rect 339 688 373 704
rect 373 688 382 704
rect 330 652 382 688
rect 486 506 538 542
rect 486 490 495 506
rect 495 490 529 506
rect 529 490 538 506
rect 486 472 495 478
rect 495 472 529 478
rect 529 472 538 478
rect 486 434 538 472
rect 486 426 495 434
rect 495 426 529 434
rect 529 426 538 434
rect 486 400 495 414
rect 495 400 529 414
rect 529 400 538 414
rect 486 362 538 400
rect 486 328 495 350
rect 495 328 529 350
rect 529 328 538 350
rect 486 298 538 328
rect 486 256 495 286
rect 495 256 529 286
rect 529 256 538 286
rect 486 234 538 256
rect 486 218 538 222
rect 486 184 495 218
rect 495 184 529 218
rect 529 184 538 218
rect 486 170 538 184
rect 486 146 538 158
rect 486 112 495 146
rect 495 112 529 146
rect 529 112 538 146
rect 486 106 538 112
rect 642 1082 694 1088
rect 642 1048 651 1082
rect 651 1048 685 1082
rect 685 1048 694 1082
rect 642 1036 694 1048
rect 642 1010 694 1024
rect 642 976 651 1010
rect 651 976 685 1010
rect 685 976 694 1010
rect 642 972 694 976
rect 642 938 694 960
rect 642 908 651 938
rect 651 908 685 938
rect 685 908 694 938
rect 642 866 694 896
rect 642 844 651 866
rect 651 844 685 866
rect 685 844 694 866
rect 642 794 694 832
rect 642 780 651 794
rect 651 780 685 794
rect 685 780 694 794
rect 642 760 651 768
rect 651 760 685 768
rect 685 760 694 768
rect 642 722 694 760
rect 642 716 651 722
rect 651 716 685 722
rect 685 716 694 722
rect 642 688 651 704
rect 651 688 685 704
rect 685 688 694 704
rect 642 652 694 688
rect 798 506 850 542
rect 798 490 807 506
rect 807 490 841 506
rect 841 490 850 506
rect 798 472 807 478
rect 807 472 841 478
rect 841 472 850 478
rect 798 434 850 472
rect 798 426 807 434
rect 807 426 841 434
rect 841 426 850 434
rect 798 400 807 414
rect 807 400 841 414
rect 841 400 850 414
rect 798 362 850 400
rect 798 328 807 350
rect 807 328 841 350
rect 841 328 850 350
rect 798 298 850 328
rect 798 256 807 286
rect 807 256 841 286
rect 841 256 850 286
rect 798 234 850 256
rect 798 218 850 222
rect 798 184 807 218
rect 807 184 841 218
rect 841 184 850 218
rect 798 170 850 184
rect 798 146 850 158
rect 798 112 807 146
rect 807 112 841 146
rect 841 112 850 146
rect 798 106 850 112
<< metal2 >>
rect 10 1088 1014 1094
rect 10 1036 330 1088
rect 382 1036 642 1088
rect 694 1036 1014 1088
rect 10 1024 1014 1036
rect 10 972 330 1024
rect 382 972 642 1024
rect 694 972 1014 1024
rect 10 960 1014 972
rect 10 908 330 960
rect 382 908 642 960
rect 694 908 1014 960
rect 10 896 1014 908
rect 10 844 330 896
rect 382 844 642 896
rect 694 844 1014 896
rect 10 832 1014 844
rect 10 780 330 832
rect 382 780 642 832
rect 694 780 1014 832
rect 10 768 1014 780
rect 10 716 330 768
rect 382 716 642 768
rect 694 716 1014 768
rect 10 704 1014 716
rect 10 652 330 704
rect 382 652 642 704
rect 694 652 1014 704
rect 10 622 1014 652
rect 10 542 1014 572
rect 10 490 174 542
rect 226 490 486 542
rect 538 490 798 542
rect 850 490 1014 542
rect 10 478 1014 490
rect 10 426 174 478
rect 226 426 486 478
rect 538 426 798 478
rect 850 426 1014 478
rect 10 414 1014 426
rect 10 362 174 414
rect 226 362 486 414
rect 538 362 798 414
rect 850 362 1014 414
rect 10 350 1014 362
rect 10 298 174 350
rect 226 298 486 350
rect 538 298 798 350
rect 850 298 1014 350
rect 10 286 1014 298
rect 10 234 174 286
rect 226 234 486 286
rect 538 234 798 286
rect 850 234 1014 286
rect 10 222 1014 234
rect 10 170 174 222
rect 226 170 486 222
rect 538 170 798 222
rect 850 170 1014 222
rect 10 158 1014 170
rect 10 106 174 158
rect 226 106 486 158
rect 538 106 798 158
rect 850 106 1014 158
rect 10 100 1014 106
<< labels >>
flabel comment s 200 597 200 597 0 FreeSans 300 0 0 0 S
flabel comment s 200 597 200 597 0 FreeSans 300 0 0 0 S
flabel comment s 356 597 356 597 0 FreeSans 300 0 0 0 S
flabel comment s 356 597 356 597 0 FreeSans 300 0 0 0 D
flabel comment s 512 597 512 597 0 FreeSans 300 0 0 0 S
flabel comment s 512 597 512 597 0 FreeSans 300 0 0 0 S
flabel comment s 668 597 668 597 0 FreeSans 300 0 0 0 S
flabel comment s 668 597 668 597 0 FreeSans 300 0 0 0 D
flabel comment s 824 597 824 597 0 FreeSans 300 0 0 0 S
flabel metal2 s 32 894 143 951 0 FreeSans 200 0 0 0 DRAIN
port 2 nsew
flabel metal2 s 32 345 134 391 0 FreeSans 200 0 0 0 SOURCE
port 3 nsew
flabel metal1 s 948 494 972 674 0 FreeSans 200 90 0 0 SUBSTRATE
port 4 nsew
flabel metal1 s 54 480 79 671 0 FreeSans 200 90 0 0 SUBSTRATE
port 4 nsew
flabel metal1 s 448 9 585 51 0 FreeSans 200 0 0 0 GATE
port 5 nsew
flabel metal1 s 443 1136 579 1176 0 FreeSans 200 0 0 0 GATE
port 5 nsew
<< properties >>
string GDS_END 7100654
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 7077692
<< end >>
