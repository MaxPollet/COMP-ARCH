magic
tech sky130A
magscale 1 2
timestamp 1681267127
<< locali >>
rect 199 732 207 766
rect 241 732 279 766
rect 313 732 351 766
rect 385 732 423 766
rect 457 732 495 766
rect 529 732 567 766
rect 601 732 639 766
rect 673 732 711 766
rect 745 732 783 766
rect 817 732 855 766
rect 889 732 927 766
rect 961 732 999 766
rect 1033 732 1071 766
rect 1105 732 1143 766
rect 1177 732 1215 766
rect 1249 732 1287 766
rect 1321 732 1359 766
rect 1393 732 1431 766
rect 1465 732 1503 766
rect 1537 732 1575 766
rect 1609 732 1647 766
rect 1681 732 1719 766
rect 1753 732 1761 766
rect 199 20 207 54
rect 241 20 279 54
rect 313 20 351 54
rect 385 20 423 54
rect 457 20 495 54
rect 529 20 567 54
rect 601 20 639 54
rect 673 20 711 54
rect 745 20 783 54
rect 817 20 855 54
rect 889 20 927 54
rect 961 20 999 54
rect 1033 20 1071 54
rect 1105 20 1143 54
rect 1177 20 1215 54
rect 1249 20 1287 54
rect 1321 20 1359 54
rect 1393 20 1431 54
rect 1465 20 1503 54
rect 1537 20 1575 54
rect 1609 20 1647 54
rect 1681 20 1719 54
rect 1753 20 1761 54
<< viali >>
rect 207 732 241 766
rect 279 732 313 766
rect 351 732 385 766
rect 423 732 457 766
rect 495 732 529 766
rect 567 732 601 766
rect 639 732 673 766
rect 711 732 745 766
rect 783 732 817 766
rect 855 732 889 766
rect 927 732 961 766
rect 999 732 1033 766
rect 1071 732 1105 766
rect 1143 732 1177 766
rect 1215 732 1249 766
rect 1287 732 1321 766
rect 1359 732 1393 766
rect 1431 732 1465 766
rect 1503 732 1537 766
rect 1575 732 1609 766
rect 1647 732 1681 766
rect 1719 732 1753 766
rect 207 20 241 54
rect 279 20 313 54
rect 351 20 385 54
rect 423 20 457 54
rect 495 20 529 54
rect 567 20 601 54
rect 639 20 673 54
rect 711 20 745 54
rect 783 20 817 54
rect 855 20 889 54
rect 927 20 961 54
rect 999 20 1033 54
rect 1071 20 1105 54
rect 1143 20 1177 54
rect 1215 20 1249 54
rect 1287 20 1321 54
rect 1359 20 1393 54
rect 1431 20 1465 54
rect 1503 20 1537 54
rect 1575 20 1609 54
rect 1647 20 1681 54
rect 1719 20 1753 54
<< obsli1 >>
rect 48 662 82 664
rect 48 590 82 628
rect 48 518 82 556
rect 48 446 82 484
rect 48 374 82 412
rect 48 302 82 340
rect 48 230 82 268
rect 48 158 82 196
rect 48 122 82 124
rect 183 88 217 698
rect 339 88 373 698
rect 495 88 529 698
rect 651 88 685 698
rect 807 88 841 698
rect 963 88 997 698
rect 1119 88 1153 698
rect 1275 88 1309 698
rect 1431 88 1465 698
rect 1587 88 1621 698
rect 1743 88 1777 698
rect 1878 662 1912 664
rect 1878 590 1912 628
rect 1878 518 1912 556
rect 1878 446 1912 484
rect 1878 374 1912 412
rect 1878 302 1912 340
rect 1878 230 1912 268
rect 1878 158 1912 196
rect 1878 122 1912 124
<< obsli1c >>
rect 48 628 82 662
rect 48 556 82 590
rect 48 484 82 518
rect 48 412 82 446
rect 48 340 82 374
rect 48 268 82 302
rect 48 196 82 230
rect 48 124 82 158
rect 1878 628 1912 662
rect 1878 556 1912 590
rect 1878 484 1912 518
rect 1878 412 1912 446
rect 1878 340 1912 374
rect 1878 268 1912 302
rect 1878 196 1912 230
rect 1878 124 1912 158
<< metal1 >>
rect 195 766 1765 786
rect 195 732 207 766
rect 241 732 279 766
rect 313 732 351 766
rect 385 732 423 766
rect 457 732 495 766
rect 529 732 567 766
rect 601 732 639 766
rect 673 732 711 766
rect 745 732 783 766
rect 817 732 855 766
rect 889 732 927 766
rect 961 732 999 766
rect 1033 732 1071 766
rect 1105 732 1143 766
rect 1177 732 1215 766
rect 1249 732 1287 766
rect 1321 732 1359 766
rect 1393 732 1431 766
rect 1465 732 1503 766
rect 1537 732 1575 766
rect 1609 732 1647 766
rect 1681 732 1719 766
rect 1753 732 1765 766
rect 195 720 1765 732
rect 36 662 94 674
rect 36 628 48 662
rect 82 628 94 662
rect 36 590 94 628
rect 36 556 48 590
rect 82 556 94 590
rect 36 518 94 556
rect 36 484 48 518
rect 82 484 94 518
rect 36 446 94 484
rect 36 412 48 446
rect 82 412 94 446
rect 36 374 94 412
rect 36 340 48 374
rect 82 340 94 374
rect 36 302 94 340
rect 36 268 48 302
rect 82 268 94 302
rect 36 230 94 268
rect 36 196 48 230
rect 82 196 94 230
rect 36 158 94 196
rect 36 124 48 158
rect 82 124 94 158
rect 36 112 94 124
rect 1866 662 1924 674
rect 1866 628 1878 662
rect 1912 628 1924 662
rect 1866 590 1924 628
rect 1866 556 1878 590
rect 1912 556 1924 590
rect 1866 518 1924 556
rect 1866 484 1878 518
rect 1912 484 1924 518
rect 1866 446 1924 484
rect 1866 412 1878 446
rect 1912 412 1924 446
rect 1866 374 1924 412
rect 1866 340 1878 374
rect 1912 340 1924 374
rect 1866 302 1924 340
rect 1866 268 1878 302
rect 1912 268 1924 302
rect 1866 230 1924 268
rect 1866 196 1878 230
rect 1912 196 1924 230
rect 1866 158 1924 196
rect 1866 124 1878 158
rect 1912 124 1924 158
rect 1866 112 1924 124
rect 195 54 1765 66
rect 195 20 207 54
rect 241 20 279 54
rect 313 20 351 54
rect 385 20 423 54
rect 457 20 495 54
rect 529 20 567 54
rect 601 20 639 54
rect 673 20 711 54
rect 745 20 783 54
rect 817 20 855 54
rect 889 20 927 54
rect 961 20 999 54
rect 1033 20 1071 54
rect 1105 20 1143 54
rect 1177 20 1215 54
rect 1249 20 1287 54
rect 1321 20 1359 54
rect 1393 20 1431 54
rect 1465 20 1503 54
rect 1537 20 1575 54
rect 1609 20 1647 54
rect 1681 20 1719 54
rect 1753 20 1765 54
rect 195 0 1765 20
<< obsm1 >>
rect 174 112 226 674
rect 330 112 382 674
rect 486 112 538 674
rect 642 112 694 674
rect 798 112 850 674
rect 954 112 1006 674
rect 1110 112 1162 674
rect 1266 112 1318 674
rect 1422 112 1474 674
rect 1578 112 1630 674
rect 1734 112 1786 674
<< metal2 >>
rect 10 418 1950 674
rect 10 112 1950 368
<< labels >>
rlabel metal2 s 10 418 1950 674 6 DRAIN
port 1 nsew
rlabel viali s 1719 732 1753 766 6 GATE
port 2 nsew
rlabel viali s 1719 20 1753 54 6 GATE
port 2 nsew
rlabel viali s 1647 732 1681 766 6 GATE
port 2 nsew
rlabel viali s 1647 20 1681 54 6 GATE
port 2 nsew
rlabel viali s 1575 732 1609 766 6 GATE
port 2 nsew
rlabel viali s 1575 20 1609 54 6 GATE
port 2 nsew
rlabel viali s 1503 732 1537 766 6 GATE
port 2 nsew
rlabel viali s 1503 20 1537 54 6 GATE
port 2 nsew
rlabel viali s 1431 732 1465 766 6 GATE
port 2 nsew
rlabel viali s 1431 20 1465 54 6 GATE
port 2 nsew
rlabel viali s 1359 732 1393 766 6 GATE
port 2 nsew
rlabel viali s 1359 20 1393 54 6 GATE
port 2 nsew
rlabel viali s 1287 732 1321 766 6 GATE
port 2 nsew
rlabel viali s 1287 20 1321 54 6 GATE
port 2 nsew
rlabel viali s 1215 732 1249 766 6 GATE
port 2 nsew
rlabel viali s 1215 20 1249 54 6 GATE
port 2 nsew
rlabel viali s 1143 732 1177 766 6 GATE
port 2 nsew
rlabel viali s 1143 20 1177 54 6 GATE
port 2 nsew
rlabel viali s 1071 732 1105 766 6 GATE
port 2 nsew
rlabel viali s 1071 20 1105 54 6 GATE
port 2 nsew
rlabel viali s 999 732 1033 766 6 GATE
port 2 nsew
rlabel viali s 999 20 1033 54 6 GATE
port 2 nsew
rlabel viali s 927 732 961 766 6 GATE
port 2 nsew
rlabel viali s 927 20 961 54 6 GATE
port 2 nsew
rlabel viali s 855 732 889 766 6 GATE
port 2 nsew
rlabel viali s 855 20 889 54 6 GATE
port 2 nsew
rlabel viali s 783 732 817 766 6 GATE
port 2 nsew
rlabel viali s 783 20 817 54 6 GATE
port 2 nsew
rlabel viali s 711 732 745 766 6 GATE
port 2 nsew
rlabel viali s 711 20 745 54 6 GATE
port 2 nsew
rlabel viali s 639 732 673 766 6 GATE
port 2 nsew
rlabel viali s 639 20 673 54 6 GATE
port 2 nsew
rlabel viali s 567 732 601 766 6 GATE
port 2 nsew
rlabel viali s 567 20 601 54 6 GATE
port 2 nsew
rlabel viali s 495 732 529 766 6 GATE
port 2 nsew
rlabel viali s 495 20 529 54 6 GATE
port 2 nsew
rlabel viali s 423 732 457 766 6 GATE
port 2 nsew
rlabel viali s 423 20 457 54 6 GATE
port 2 nsew
rlabel viali s 351 732 385 766 6 GATE
port 2 nsew
rlabel viali s 351 20 385 54 6 GATE
port 2 nsew
rlabel viali s 279 732 313 766 6 GATE
port 2 nsew
rlabel viali s 279 20 313 54 6 GATE
port 2 nsew
rlabel viali s 207 732 241 766 6 GATE
port 2 nsew
rlabel viali s 207 20 241 54 6 GATE
port 2 nsew
rlabel locali s 199 732 1761 766 6 GATE
port 2 nsew
rlabel locali s 199 20 1761 54 6 GATE
port 2 nsew
rlabel metal1 s 195 720 1765 786 6 GATE
port 2 nsew
rlabel metal1 s 195 0 1765 66 6 GATE
port 2 nsew
rlabel metal2 s 10 112 1950 368 6 SOURCE
port 3 nsew
rlabel metal1 s 36 112 94 674 6 SUBSTRATE
port 4 nsew
rlabel metal1 s 1866 112 1924 674 6 SUBSTRATE
port 4 nsew
<< properties >>
string FIXED_BBOX 10 0 1950 786
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 7776296
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 7744842
<< end >>
