magic
tech sky130A
magscale 1 2
timestamp 1681267127
<< nwell >>
rect -38 261 2430 582
<< pwell >>
rect 1924 201 2391 203
rect 782 157 1236 201
rect 1557 157 2391 201
rect 1 21 2391 157
rect 30 -17 64 21
<< locali >>
rect 17 195 88 325
rect 350 201 432 325
rect 2040 326 2097 493
rect 1863 219 1938 265
rect 2056 143 2097 326
rect 2040 51 2097 143
rect 2323 289 2375 493
rect 2332 165 2375 289
rect 2323 51 2375 165
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2392 561
rect 17 393 69 493
rect 103 427 169 527
rect 17 359 168 393
rect 122 161 168 359
rect 17 127 168 161
rect 17 69 69 127
rect 103 17 169 93
rect 203 69 248 493
rect 287 427 357 527
rect 391 393 425 493
rect 468 450 634 484
rect 282 359 425 393
rect 282 165 316 359
rect 466 315 566 391
rect 282 127 425 165
rect 466 141 510 315
rect 600 281 634 450
rect 682 441 758 527
rect 818 407 852 475
rect 668 357 938 407
rect 976 383 1042 527
rect 1251 450 1417 484
rect 1465 451 1541 527
rect 668 315 718 357
rect 820 281 870 297
rect 600 247 870 281
rect 600 239 680 247
rect 546 129 612 203
rect 287 17 357 93
rect 391 61 425 127
rect 646 93 680 239
rect 826 231 870 247
rect 904 213 938 357
rect 972 283 1173 331
rect 1213 315 1260 397
rect 972 247 1038 283
rect 1308 261 1349 381
rect 1100 213 1166 247
rect 718 193 784 213
rect 718 187 800 193
rect 718 153 766 187
rect 904 179 1166 213
rect 1225 225 1349 261
rect 1383 281 1417 450
rect 1589 417 1623 475
rect 1729 451 2006 527
rect 1451 383 2006 417
rect 1451 315 1501 383
rect 1383 247 1653 281
rect 904 153 948 179
rect 718 147 800 153
rect 882 119 948 153
rect 481 53 680 93
rect 714 17 748 105
rect 782 85 848 109
rect 982 85 1016 143
rect 1225 141 1282 225
rect 1383 93 1417 247
rect 1609 215 1653 247
rect 1492 187 1567 213
rect 1492 153 1502 187
rect 1536 153 1567 187
rect 1687 156 1723 383
rect 1492 147 1567 153
rect 1657 119 1723 156
rect 1757 315 1909 349
rect 1757 185 1812 315
rect 1972 265 2006 383
rect 1972 199 2022 265
rect 1757 151 1895 185
rect 782 51 1016 85
rect 1070 17 1136 93
rect 1264 53 1417 93
rect 1453 17 1505 105
rect 1557 85 1623 109
rect 1757 85 1791 117
rect 1557 51 1791 85
rect 1848 53 1895 151
rect 1940 17 2006 161
rect 2131 265 2194 483
rect 2230 353 2289 527
rect 2131 199 2298 265
rect 2131 51 2194 199
rect 2230 17 2289 109
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2392 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 766 153 800 187
rect 1502 153 1536 187
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
<< metal1 >>
rect 0 561 2392 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2392 561
rect 0 496 2392 527
rect 754 187 812 193
rect 754 153 766 187
rect 800 184 812 187
rect 1490 187 1548 193
rect 1490 184 1502 187
rect 800 156 1502 184
rect 800 153 812 156
rect 754 147 812 153
rect 1490 153 1502 156
rect 1536 153 1548 187
rect 1490 147 1548 153
rect 0 17 2392 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2392 17
rect 0 -48 2392 -17
<< obsm1 >>
rect 110 388 168 397
rect 478 388 536 397
rect 1214 388 1272 397
rect 110 360 1272 388
rect 110 351 168 360
rect 478 351 536 360
rect 1214 351 1272 360
rect 1122 320 1180 329
rect 1766 320 1824 329
rect 1122 292 1824 320
rect 1122 283 1180 292
rect 1766 283 1824 292
rect 1214 252 1272 261
rect 585 224 1272 252
rect 585 193 624 224
rect 1214 215 1272 224
rect 202 184 260 193
rect 566 184 624 193
rect 202 156 624 184
rect 202 147 260 156
rect 566 147 624 156
<< labels >>
rlabel locali s 17 195 88 325 6 CLK
port 1 nsew clock input
rlabel locali s 350 201 432 325 6 D
port 2 nsew signal input
rlabel locali s 1863 219 1938 265 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 1490 147 1548 156 6 SET_B
port 4 nsew signal input
rlabel metal1 s 754 147 812 156 6 SET_B
port 4 nsew signal input
rlabel metal1 s 754 156 1548 184 6 SET_B
port 4 nsew signal input
rlabel metal1 s 1490 184 1548 193 6 SET_B
port 4 nsew signal input
rlabel metal1 s 754 184 812 193 6 SET_B
port 4 nsew signal input
rlabel metal1 s 0 -48 2392 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1 21 2391 157 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1557 157 2391 201 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 782 157 1236 201 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1924 201 2391 203 6 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 2430 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 2392 592 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 2323 51 2375 165 6 Q
port 9 nsew signal output
rlabel locali s 2332 165 2375 289 6 Q
port 9 nsew signal output
rlabel locali s 2323 289 2375 493 6 Q
port 9 nsew signal output
rlabel locali s 2040 51 2097 143 6 Q_N
port 10 nsew signal output
rlabel locali s 2056 143 2097 326 6 Q_N
port 10 nsew signal output
rlabel locali s 2040 326 2097 493 6 Q_N
port 10 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 2392 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 3423836
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3404818
<< end >>
