magic
tech sky130A
magscale 1 2
timestamp 1681267127
use sky130_fd_pr__hvdfl1sd2__example_55959141808306  sky130_fd_pr__hvdfl1sd2__example_55959141808306_0
timestamp 1681267127
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808306  sky130_fd_pr__hvdfl1sd2__example_55959141808306_1
timestamp 1681267127
transform 1 0 100 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 8081174
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 8080244
<< end >>
