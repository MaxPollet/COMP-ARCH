magic
tech sky130A
timestamp 1681267127
<< properties >>
string GDS_END 38343208
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 38342504
<< end >>
