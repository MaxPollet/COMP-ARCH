magic
tech sky130A
magscale 1 2
timestamp 1681267127
<< nwell >>
rect 415 600 14720 4720
<< pwell >>
rect 10 4857 15126 5109
rect 10 540 355 4857
rect 14781 540 15126 4857
rect 10 288 15126 540
<< mvpmos >>
rect 881 3152 1001 4152
rect 1311 3152 1431 4152
rect 1873 3152 1993 4152
rect 2303 3152 2423 4152
rect 2865 3152 2985 4152
rect 3295 3152 3415 4152
rect 3857 3152 3977 4152
rect 4287 3152 4407 4152
rect 4849 3152 4969 4152
rect 5279 3152 5399 4152
rect 5841 3152 5961 4152
rect 6271 3152 6391 4152
rect 6833 3152 6953 4152
rect 7263 3152 7383 4152
rect 7825 3152 7945 4152
rect 8255 3152 8375 4152
rect 8817 3152 8937 4152
rect 9247 3152 9367 4152
rect 9809 3152 9929 4152
rect 10239 3152 10359 4152
rect 10801 3152 10921 4152
rect 11231 3152 11351 4152
rect 11793 3152 11913 4152
rect 12223 3152 12343 4152
rect 12785 3152 12905 4152
rect 13215 3152 13335 4152
rect 13777 3152 13897 4152
rect 14135 3152 14255 4152
rect 881 1552 1001 2552
rect 1311 1552 1431 2552
rect 1873 1552 1993 2552
rect 2303 1552 2423 2552
rect 2865 1552 2985 2552
rect 3295 1552 3415 2552
rect 3857 1552 3977 2552
rect 4287 1552 4407 2552
rect 4849 1552 4969 2552
rect 5279 1552 5399 2552
rect 5841 1552 5961 2552
rect 6271 1552 6391 2552
rect 6833 1552 6953 2552
rect 7263 1552 7383 2552
rect 7825 1552 7945 2552
rect 8255 1552 8375 2552
rect 8817 1552 8937 2552
rect 9247 1552 9367 2552
rect 9809 1552 9929 2552
rect 10239 1552 10359 2552
rect 10801 1552 10921 2552
rect 11231 1552 11351 2552
rect 11793 1552 11913 2552
rect 12223 1552 12343 2552
rect 12785 1552 12905 2552
rect 13215 1552 13335 2552
rect 13777 1552 13897 2552
rect 14135 1552 14255 2552
<< mvpdiff >>
rect 708 4082 881 4152
rect 708 4048 745 4082
rect 779 4048 881 4082
rect 708 4014 881 4048
rect 708 3980 745 4014
rect 779 3980 881 4014
rect 708 3946 881 3980
rect 708 3912 745 3946
rect 779 3912 881 3946
rect 708 3878 881 3912
rect 708 3844 745 3878
rect 779 3844 881 3878
rect 708 3810 881 3844
rect 708 3776 745 3810
rect 779 3776 881 3810
rect 708 3742 881 3776
rect 708 3708 745 3742
rect 779 3708 881 3742
rect 708 3674 881 3708
rect 708 3640 745 3674
rect 779 3640 881 3674
rect 708 3606 881 3640
rect 708 3572 745 3606
rect 779 3572 881 3606
rect 708 3538 881 3572
rect 708 3504 745 3538
rect 779 3504 881 3538
rect 708 3470 881 3504
rect 708 3436 745 3470
rect 779 3436 881 3470
rect 708 3402 881 3436
rect 708 3368 745 3402
rect 779 3368 881 3402
rect 708 3334 881 3368
rect 708 3300 745 3334
rect 779 3300 881 3334
rect 708 3266 881 3300
rect 708 3232 745 3266
rect 779 3232 881 3266
rect 708 3198 881 3232
rect 708 3164 745 3198
rect 779 3164 881 3198
rect 708 3152 881 3164
rect 1001 4082 1311 4152
rect 1001 4048 1103 4082
rect 1137 4048 1175 4082
rect 1209 4048 1311 4082
rect 1001 4014 1311 4048
rect 1001 3980 1103 4014
rect 1137 3980 1175 4014
rect 1209 3980 1311 4014
rect 1001 3946 1311 3980
rect 1001 3912 1103 3946
rect 1137 3912 1175 3946
rect 1209 3912 1311 3946
rect 1001 3878 1311 3912
rect 1001 3844 1103 3878
rect 1137 3844 1175 3878
rect 1209 3844 1311 3878
rect 1001 3810 1311 3844
rect 1001 3776 1103 3810
rect 1137 3776 1175 3810
rect 1209 3776 1311 3810
rect 1001 3742 1311 3776
rect 1001 3708 1103 3742
rect 1137 3708 1175 3742
rect 1209 3708 1311 3742
rect 1001 3674 1311 3708
rect 1001 3640 1103 3674
rect 1137 3640 1175 3674
rect 1209 3640 1311 3674
rect 1001 3606 1311 3640
rect 1001 3572 1103 3606
rect 1137 3572 1175 3606
rect 1209 3572 1311 3606
rect 1001 3538 1311 3572
rect 1001 3504 1103 3538
rect 1137 3504 1175 3538
rect 1209 3504 1311 3538
rect 1001 3470 1311 3504
rect 1001 3436 1103 3470
rect 1137 3436 1175 3470
rect 1209 3436 1311 3470
rect 1001 3402 1311 3436
rect 1001 3368 1103 3402
rect 1137 3368 1175 3402
rect 1209 3368 1311 3402
rect 1001 3334 1311 3368
rect 1001 3300 1103 3334
rect 1137 3300 1175 3334
rect 1209 3300 1311 3334
rect 1001 3266 1311 3300
rect 1001 3232 1103 3266
rect 1137 3232 1175 3266
rect 1209 3232 1311 3266
rect 1001 3198 1311 3232
rect 1001 3164 1103 3198
rect 1137 3164 1175 3198
rect 1209 3164 1311 3198
rect 1001 3152 1311 3164
rect 1431 4082 1582 4152
rect 1722 4082 1873 4152
rect 1431 4048 1533 4082
rect 1567 4048 1582 4082
rect 1722 4048 1737 4082
rect 1771 4048 1873 4082
rect 1431 4014 1582 4048
rect 1722 4014 1873 4048
rect 1431 3980 1533 4014
rect 1567 3980 1582 4014
rect 1722 3980 1737 4014
rect 1771 3980 1873 4014
rect 1431 3946 1582 3980
rect 1722 3946 1873 3980
rect 1431 3912 1533 3946
rect 1567 3912 1582 3946
rect 1722 3912 1737 3946
rect 1771 3912 1873 3946
rect 1431 3878 1582 3912
rect 1722 3878 1873 3912
rect 1431 3844 1533 3878
rect 1567 3844 1582 3878
rect 1722 3844 1737 3878
rect 1771 3844 1873 3878
rect 1431 3810 1582 3844
rect 1722 3810 1873 3844
rect 1431 3776 1533 3810
rect 1567 3776 1582 3810
rect 1722 3776 1737 3810
rect 1771 3776 1873 3810
rect 1431 3742 1582 3776
rect 1722 3742 1873 3776
rect 1431 3708 1533 3742
rect 1567 3708 1582 3742
rect 1722 3708 1737 3742
rect 1771 3708 1873 3742
rect 1431 3674 1582 3708
rect 1722 3674 1873 3708
rect 1431 3640 1533 3674
rect 1567 3640 1582 3674
rect 1722 3640 1737 3674
rect 1771 3640 1873 3674
rect 1431 3606 1582 3640
rect 1722 3606 1873 3640
rect 1431 3572 1533 3606
rect 1567 3572 1582 3606
rect 1722 3572 1737 3606
rect 1771 3572 1873 3606
rect 1431 3538 1582 3572
rect 1722 3538 1873 3572
rect 1431 3504 1533 3538
rect 1567 3504 1582 3538
rect 1722 3504 1737 3538
rect 1771 3504 1873 3538
rect 1431 3470 1582 3504
rect 1722 3470 1873 3504
rect 1431 3436 1533 3470
rect 1567 3436 1582 3470
rect 1722 3436 1737 3470
rect 1771 3436 1873 3470
rect 1431 3402 1582 3436
rect 1722 3402 1873 3436
rect 1431 3368 1533 3402
rect 1567 3368 1582 3402
rect 1722 3368 1737 3402
rect 1771 3368 1873 3402
rect 1431 3334 1582 3368
rect 1722 3334 1873 3368
rect 1431 3300 1533 3334
rect 1567 3300 1582 3334
rect 1722 3300 1737 3334
rect 1771 3300 1873 3334
rect 1431 3266 1582 3300
rect 1722 3266 1873 3300
rect 1431 3232 1533 3266
rect 1567 3232 1582 3266
rect 1722 3232 1737 3266
rect 1771 3232 1873 3266
rect 1431 3198 1582 3232
rect 1722 3198 1873 3232
rect 1431 3164 1533 3198
rect 1567 3164 1582 3198
rect 1722 3164 1737 3198
rect 1771 3164 1873 3198
rect 1431 3152 1582 3164
rect 1722 3152 1873 3164
rect 1993 4082 2303 4152
rect 1993 4048 2095 4082
rect 2129 4048 2167 4082
rect 2201 4048 2303 4082
rect 1993 4014 2303 4048
rect 1993 3980 2095 4014
rect 2129 3980 2167 4014
rect 2201 3980 2303 4014
rect 1993 3946 2303 3980
rect 1993 3912 2095 3946
rect 2129 3912 2167 3946
rect 2201 3912 2303 3946
rect 1993 3878 2303 3912
rect 1993 3844 2095 3878
rect 2129 3844 2167 3878
rect 2201 3844 2303 3878
rect 1993 3810 2303 3844
rect 1993 3776 2095 3810
rect 2129 3776 2167 3810
rect 2201 3776 2303 3810
rect 1993 3742 2303 3776
rect 1993 3708 2095 3742
rect 2129 3708 2167 3742
rect 2201 3708 2303 3742
rect 1993 3674 2303 3708
rect 1993 3640 2095 3674
rect 2129 3640 2167 3674
rect 2201 3640 2303 3674
rect 1993 3606 2303 3640
rect 1993 3572 2095 3606
rect 2129 3572 2167 3606
rect 2201 3572 2303 3606
rect 1993 3538 2303 3572
rect 1993 3504 2095 3538
rect 2129 3504 2167 3538
rect 2201 3504 2303 3538
rect 1993 3470 2303 3504
rect 1993 3436 2095 3470
rect 2129 3436 2167 3470
rect 2201 3436 2303 3470
rect 1993 3402 2303 3436
rect 1993 3368 2095 3402
rect 2129 3368 2167 3402
rect 2201 3368 2303 3402
rect 1993 3334 2303 3368
rect 1993 3300 2095 3334
rect 2129 3300 2167 3334
rect 2201 3300 2303 3334
rect 1993 3266 2303 3300
rect 1993 3232 2095 3266
rect 2129 3232 2167 3266
rect 2201 3232 2303 3266
rect 1993 3198 2303 3232
rect 1993 3164 2095 3198
rect 2129 3164 2167 3198
rect 2201 3164 2303 3198
rect 1993 3152 2303 3164
rect 2423 4082 2574 4152
rect 2714 4082 2865 4152
rect 2423 4048 2525 4082
rect 2559 4048 2574 4082
rect 2714 4048 2729 4082
rect 2763 4048 2865 4082
rect 2423 4014 2574 4048
rect 2714 4014 2865 4048
rect 2423 3980 2525 4014
rect 2559 3980 2574 4014
rect 2714 3980 2729 4014
rect 2763 3980 2865 4014
rect 2423 3946 2574 3980
rect 2714 3946 2865 3980
rect 2423 3912 2525 3946
rect 2559 3912 2574 3946
rect 2714 3912 2729 3946
rect 2763 3912 2865 3946
rect 2423 3878 2574 3912
rect 2714 3878 2865 3912
rect 2423 3844 2525 3878
rect 2559 3844 2574 3878
rect 2714 3844 2729 3878
rect 2763 3844 2865 3878
rect 2423 3810 2574 3844
rect 2714 3810 2865 3844
rect 2423 3776 2525 3810
rect 2559 3776 2574 3810
rect 2714 3776 2729 3810
rect 2763 3776 2865 3810
rect 2423 3742 2574 3776
rect 2714 3742 2865 3776
rect 2423 3708 2525 3742
rect 2559 3708 2574 3742
rect 2714 3708 2729 3742
rect 2763 3708 2865 3742
rect 2423 3674 2574 3708
rect 2714 3674 2865 3708
rect 2423 3640 2525 3674
rect 2559 3640 2574 3674
rect 2714 3640 2729 3674
rect 2763 3640 2865 3674
rect 2423 3606 2574 3640
rect 2714 3606 2865 3640
rect 2423 3572 2525 3606
rect 2559 3572 2574 3606
rect 2714 3572 2729 3606
rect 2763 3572 2865 3606
rect 2423 3538 2574 3572
rect 2714 3538 2865 3572
rect 2423 3504 2525 3538
rect 2559 3504 2574 3538
rect 2714 3504 2729 3538
rect 2763 3504 2865 3538
rect 2423 3470 2574 3504
rect 2714 3470 2865 3504
rect 2423 3436 2525 3470
rect 2559 3436 2574 3470
rect 2714 3436 2729 3470
rect 2763 3436 2865 3470
rect 2423 3402 2574 3436
rect 2714 3402 2865 3436
rect 2423 3368 2525 3402
rect 2559 3368 2574 3402
rect 2714 3368 2729 3402
rect 2763 3368 2865 3402
rect 2423 3334 2574 3368
rect 2714 3334 2865 3368
rect 2423 3300 2525 3334
rect 2559 3300 2574 3334
rect 2714 3300 2729 3334
rect 2763 3300 2865 3334
rect 2423 3266 2574 3300
rect 2714 3266 2865 3300
rect 2423 3232 2525 3266
rect 2559 3232 2574 3266
rect 2714 3232 2729 3266
rect 2763 3232 2865 3266
rect 2423 3198 2574 3232
rect 2714 3198 2865 3232
rect 2423 3164 2525 3198
rect 2559 3164 2574 3198
rect 2714 3164 2729 3198
rect 2763 3164 2865 3198
rect 2423 3152 2574 3164
rect 2714 3152 2865 3164
rect 2985 4082 3295 4152
rect 2985 4048 3087 4082
rect 3121 4048 3159 4082
rect 3193 4048 3295 4082
rect 2985 4014 3295 4048
rect 2985 3980 3087 4014
rect 3121 3980 3159 4014
rect 3193 3980 3295 4014
rect 2985 3946 3295 3980
rect 2985 3912 3087 3946
rect 3121 3912 3159 3946
rect 3193 3912 3295 3946
rect 2985 3878 3295 3912
rect 2985 3844 3087 3878
rect 3121 3844 3159 3878
rect 3193 3844 3295 3878
rect 2985 3810 3295 3844
rect 2985 3776 3087 3810
rect 3121 3776 3159 3810
rect 3193 3776 3295 3810
rect 2985 3742 3295 3776
rect 2985 3708 3087 3742
rect 3121 3708 3159 3742
rect 3193 3708 3295 3742
rect 2985 3674 3295 3708
rect 2985 3640 3087 3674
rect 3121 3640 3159 3674
rect 3193 3640 3295 3674
rect 2985 3606 3295 3640
rect 2985 3572 3087 3606
rect 3121 3572 3159 3606
rect 3193 3572 3295 3606
rect 2985 3538 3295 3572
rect 2985 3504 3087 3538
rect 3121 3504 3159 3538
rect 3193 3504 3295 3538
rect 2985 3470 3295 3504
rect 2985 3436 3087 3470
rect 3121 3436 3159 3470
rect 3193 3436 3295 3470
rect 2985 3402 3295 3436
rect 2985 3368 3087 3402
rect 3121 3368 3159 3402
rect 3193 3368 3295 3402
rect 2985 3334 3295 3368
rect 2985 3300 3087 3334
rect 3121 3300 3159 3334
rect 3193 3300 3295 3334
rect 2985 3266 3295 3300
rect 2985 3232 3087 3266
rect 3121 3232 3159 3266
rect 3193 3232 3295 3266
rect 2985 3198 3295 3232
rect 2985 3164 3087 3198
rect 3121 3164 3159 3198
rect 3193 3164 3295 3198
rect 2985 3152 3295 3164
rect 3415 4082 3566 4152
rect 3706 4082 3857 4152
rect 3415 4048 3517 4082
rect 3551 4048 3566 4082
rect 3706 4048 3721 4082
rect 3755 4048 3857 4082
rect 3415 4014 3566 4048
rect 3706 4014 3857 4048
rect 3415 3980 3517 4014
rect 3551 3980 3566 4014
rect 3706 3980 3721 4014
rect 3755 3980 3857 4014
rect 3415 3946 3566 3980
rect 3706 3946 3857 3980
rect 3415 3912 3517 3946
rect 3551 3912 3566 3946
rect 3706 3912 3721 3946
rect 3755 3912 3857 3946
rect 3415 3878 3566 3912
rect 3706 3878 3857 3912
rect 3415 3844 3517 3878
rect 3551 3844 3566 3878
rect 3706 3844 3721 3878
rect 3755 3844 3857 3878
rect 3415 3810 3566 3844
rect 3706 3810 3857 3844
rect 3415 3776 3517 3810
rect 3551 3776 3566 3810
rect 3706 3776 3721 3810
rect 3755 3776 3857 3810
rect 3415 3742 3566 3776
rect 3706 3742 3857 3776
rect 3415 3708 3517 3742
rect 3551 3708 3566 3742
rect 3706 3708 3721 3742
rect 3755 3708 3857 3742
rect 3415 3674 3566 3708
rect 3706 3674 3857 3708
rect 3415 3640 3517 3674
rect 3551 3640 3566 3674
rect 3706 3640 3721 3674
rect 3755 3640 3857 3674
rect 3415 3606 3566 3640
rect 3706 3606 3857 3640
rect 3415 3572 3517 3606
rect 3551 3572 3566 3606
rect 3706 3572 3721 3606
rect 3755 3572 3857 3606
rect 3415 3538 3566 3572
rect 3706 3538 3857 3572
rect 3415 3504 3517 3538
rect 3551 3504 3566 3538
rect 3706 3504 3721 3538
rect 3755 3504 3857 3538
rect 3415 3470 3566 3504
rect 3706 3470 3857 3504
rect 3415 3436 3517 3470
rect 3551 3436 3566 3470
rect 3706 3436 3721 3470
rect 3755 3436 3857 3470
rect 3415 3402 3566 3436
rect 3706 3402 3857 3436
rect 3415 3368 3517 3402
rect 3551 3368 3566 3402
rect 3706 3368 3721 3402
rect 3755 3368 3857 3402
rect 3415 3334 3566 3368
rect 3706 3334 3857 3368
rect 3415 3300 3517 3334
rect 3551 3300 3566 3334
rect 3706 3300 3721 3334
rect 3755 3300 3857 3334
rect 3415 3266 3566 3300
rect 3706 3266 3857 3300
rect 3415 3232 3517 3266
rect 3551 3232 3566 3266
rect 3706 3232 3721 3266
rect 3755 3232 3857 3266
rect 3415 3198 3566 3232
rect 3706 3198 3857 3232
rect 3415 3164 3517 3198
rect 3551 3164 3566 3198
rect 3706 3164 3721 3198
rect 3755 3164 3857 3198
rect 3415 3152 3566 3164
rect 3706 3152 3857 3164
rect 3977 4082 4287 4152
rect 3977 4048 4079 4082
rect 4113 4048 4151 4082
rect 4185 4048 4287 4082
rect 3977 4014 4287 4048
rect 3977 3980 4079 4014
rect 4113 3980 4151 4014
rect 4185 3980 4287 4014
rect 3977 3946 4287 3980
rect 3977 3912 4079 3946
rect 4113 3912 4151 3946
rect 4185 3912 4287 3946
rect 3977 3878 4287 3912
rect 3977 3844 4079 3878
rect 4113 3844 4151 3878
rect 4185 3844 4287 3878
rect 3977 3810 4287 3844
rect 3977 3776 4079 3810
rect 4113 3776 4151 3810
rect 4185 3776 4287 3810
rect 3977 3742 4287 3776
rect 3977 3708 4079 3742
rect 4113 3708 4151 3742
rect 4185 3708 4287 3742
rect 3977 3674 4287 3708
rect 3977 3640 4079 3674
rect 4113 3640 4151 3674
rect 4185 3640 4287 3674
rect 3977 3606 4287 3640
rect 3977 3572 4079 3606
rect 4113 3572 4151 3606
rect 4185 3572 4287 3606
rect 3977 3538 4287 3572
rect 3977 3504 4079 3538
rect 4113 3504 4151 3538
rect 4185 3504 4287 3538
rect 3977 3470 4287 3504
rect 3977 3436 4079 3470
rect 4113 3436 4151 3470
rect 4185 3436 4287 3470
rect 3977 3402 4287 3436
rect 3977 3368 4079 3402
rect 4113 3368 4151 3402
rect 4185 3368 4287 3402
rect 3977 3334 4287 3368
rect 3977 3300 4079 3334
rect 4113 3300 4151 3334
rect 4185 3300 4287 3334
rect 3977 3266 4287 3300
rect 3977 3232 4079 3266
rect 4113 3232 4151 3266
rect 4185 3232 4287 3266
rect 3977 3198 4287 3232
rect 3977 3164 4079 3198
rect 4113 3164 4151 3198
rect 4185 3164 4287 3198
rect 3977 3152 4287 3164
rect 4407 4082 4558 4152
rect 4698 4082 4849 4152
rect 4407 4048 4509 4082
rect 4543 4048 4558 4082
rect 4698 4048 4713 4082
rect 4747 4048 4849 4082
rect 4407 4014 4558 4048
rect 4698 4014 4849 4048
rect 4407 3980 4509 4014
rect 4543 3980 4558 4014
rect 4698 3980 4713 4014
rect 4747 3980 4849 4014
rect 4407 3946 4558 3980
rect 4698 3946 4849 3980
rect 4407 3912 4509 3946
rect 4543 3912 4558 3946
rect 4698 3912 4713 3946
rect 4747 3912 4849 3946
rect 4407 3878 4558 3912
rect 4698 3878 4849 3912
rect 4407 3844 4509 3878
rect 4543 3844 4558 3878
rect 4698 3844 4713 3878
rect 4747 3844 4849 3878
rect 4407 3810 4558 3844
rect 4698 3810 4849 3844
rect 4407 3776 4509 3810
rect 4543 3776 4558 3810
rect 4698 3776 4713 3810
rect 4747 3776 4849 3810
rect 4407 3742 4558 3776
rect 4698 3742 4849 3776
rect 4407 3708 4509 3742
rect 4543 3708 4558 3742
rect 4698 3708 4713 3742
rect 4747 3708 4849 3742
rect 4407 3674 4558 3708
rect 4698 3674 4849 3708
rect 4407 3640 4509 3674
rect 4543 3640 4558 3674
rect 4698 3640 4713 3674
rect 4747 3640 4849 3674
rect 4407 3606 4558 3640
rect 4698 3606 4849 3640
rect 4407 3572 4509 3606
rect 4543 3572 4558 3606
rect 4698 3572 4713 3606
rect 4747 3572 4849 3606
rect 4407 3538 4558 3572
rect 4698 3538 4849 3572
rect 4407 3504 4509 3538
rect 4543 3504 4558 3538
rect 4698 3504 4713 3538
rect 4747 3504 4849 3538
rect 4407 3470 4558 3504
rect 4698 3470 4849 3504
rect 4407 3436 4509 3470
rect 4543 3436 4558 3470
rect 4698 3436 4713 3470
rect 4747 3436 4849 3470
rect 4407 3402 4558 3436
rect 4698 3402 4849 3436
rect 4407 3368 4509 3402
rect 4543 3368 4558 3402
rect 4698 3368 4713 3402
rect 4747 3368 4849 3402
rect 4407 3334 4558 3368
rect 4698 3334 4849 3368
rect 4407 3300 4509 3334
rect 4543 3300 4558 3334
rect 4698 3300 4713 3334
rect 4747 3300 4849 3334
rect 4407 3266 4558 3300
rect 4698 3266 4849 3300
rect 4407 3232 4509 3266
rect 4543 3232 4558 3266
rect 4698 3232 4713 3266
rect 4747 3232 4849 3266
rect 4407 3198 4558 3232
rect 4698 3198 4849 3232
rect 4407 3164 4509 3198
rect 4543 3164 4558 3198
rect 4698 3164 4713 3198
rect 4747 3164 4849 3198
rect 4407 3152 4558 3164
rect 4698 3152 4849 3164
rect 4969 4082 5279 4152
rect 4969 4048 5071 4082
rect 5105 4048 5143 4082
rect 5177 4048 5279 4082
rect 4969 4014 5279 4048
rect 4969 3980 5071 4014
rect 5105 3980 5143 4014
rect 5177 3980 5279 4014
rect 4969 3946 5279 3980
rect 4969 3912 5071 3946
rect 5105 3912 5143 3946
rect 5177 3912 5279 3946
rect 4969 3878 5279 3912
rect 4969 3844 5071 3878
rect 5105 3844 5143 3878
rect 5177 3844 5279 3878
rect 4969 3810 5279 3844
rect 4969 3776 5071 3810
rect 5105 3776 5143 3810
rect 5177 3776 5279 3810
rect 4969 3742 5279 3776
rect 4969 3708 5071 3742
rect 5105 3708 5143 3742
rect 5177 3708 5279 3742
rect 4969 3674 5279 3708
rect 4969 3640 5071 3674
rect 5105 3640 5143 3674
rect 5177 3640 5279 3674
rect 4969 3606 5279 3640
rect 4969 3572 5071 3606
rect 5105 3572 5143 3606
rect 5177 3572 5279 3606
rect 4969 3538 5279 3572
rect 4969 3504 5071 3538
rect 5105 3504 5143 3538
rect 5177 3504 5279 3538
rect 4969 3470 5279 3504
rect 4969 3436 5071 3470
rect 5105 3436 5143 3470
rect 5177 3436 5279 3470
rect 4969 3402 5279 3436
rect 4969 3368 5071 3402
rect 5105 3368 5143 3402
rect 5177 3368 5279 3402
rect 4969 3334 5279 3368
rect 4969 3300 5071 3334
rect 5105 3300 5143 3334
rect 5177 3300 5279 3334
rect 4969 3266 5279 3300
rect 4969 3232 5071 3266
rect 5105 3232 5143 3266
rect 5177 3232 5279 3266
rect 4969 3198 5279 3232
rect 4969 3164 5071 3198
rect 5105 3164 5143 3198
rect 5177 3164 5279 3198
rect 4969 3152 5279 3164
rect 5399 4082 5550 4152
rect 5690 4082 5841 4152
rect 5399 4048 5501 4082
rect 5535 4048 5550 4082
rect 5690 4048 5705 4082
rect 5739 4048 5841 4082
rect 5399 4014 5550 4048
rect 5690 4014 5841 4048
rect 5399 3980 5501 4014
rect 5535 3980 5550 4014
rect 5690 3980 5705 4014
rect 5739 3980 5841 4014
rect 5399 3946 5550 3980
rect 5690 3946 5841 3980
rect 5399 3912 5501 3946
rect 5535 3912 5550 3946
rect 5690 3912 5705 3946
rect 5739 3912 5841 3946
rect 5399 3878 5550 3912
rect 5690 3878 5841 3912
rect 5399 3844 5501 3878
rect 5535 3844 5550 3878
rect 5690 3844 5705 3878
rect 5739 3844 5841 3878
rect 5399 3810 5550 3844
rect 5690 3810 5841 3844
rect 5399 3776 5501 3810
rect 5535 3776 5550 3810
rect 5690 3776 5705 3810
rect 5739 3776 5841 3810
rect 5399 3742 5550 3776
rect 5690 3742 5841 3776
rect 5399 3708 5501 3742
rect 5535 3708 5550 3742
rect 5690 3708 5705 3742
rect 5739 3708 5841 3742
rect 5399 3674 5550 3708
rect 5690 3674 5841 3708
rect 5399 3640 5501 3674
rect 5535 3640 5550 3674
rect 5690 3640 5705 3674
rect 5739 3640 5841 3674
rect 5399 3606 5550 3640
rect 5690 3606 5841 3640
rect 5399 3572 5501 3606
rect 5535 3572 5550 3606
rect 5690 3572 5705 3606
rect 5739 3572 5841 3606
rect 5399 3538 5550 3572
rect 5690 3538 5841 3572
rect 5399 3504 5501 3538
rect 5535 3504 5550 3538
rect 5690 3504 5705 3538
rect 5739 3504 5841 3538
rect 5399 3470 5550 3504
rect 5690 3470 5841 3504
rect 5399 3436 5501 3470
rect 5535 3436 5550 3470
rect 5690 3436 5705 3470
rect 5739 3436 5841 3470
rect 5399 3402 5550 3436
rect 5690 3402 5841 3436
rect 5399 3368 5501 3402
rect 5535 3368 5550 3402
rect 5690 3368 5705 3402
rect 5739 3368 5841 3402
rect 5399 3334 5550 3368
rect 5690 3334 5841 3368
rect 5399 3300 5501 3334
rect 5535 3300 5550 3334
rect 5690 3300 5705 3334
rect 5739 3300 5841 3334
rect 5399 3266 5550 3300
rect 5690 3266 5841 3300
rect 5399 3232 5501 3266
rect 5535 3232 5550 3266
rect 5690 3232 5705 3266
rect 5739 3232 5841 3266
rect 5399 3198 5550 3232
rect 5690 3198 5841 3232
rect 5399 3164 5501 3198
rect 5535 3164 5550 3198
rect 5690 3164 5705 3198
rect 5739 3164 5841 3198
rect 5399 3152 5550 3164
rect 5690 3152 5841 3164
rect 5961 4082 6271 4152
rect 5961 4048 6063 4082
rect 6097 4048 6135 4082
rect 6169 4048 6271 4082
rect 5961 4014 6271 4048
rect 5961 3980 6063 4014
rect 6097 3980 6135 4014
rect 6169 3980 6271 4014
rect 5961 3946 6271 3980
rect 5961 3912 6063 3946
rect 6097 3912 6135 3946
rect 6169 3912 6271 3946
rect 5961 3878 6271 3912
rect 5961 3844 6063 3878
rect 6097 3844 6135 3878
rect 6169 3844 6271 3878
rect 5961 3810 6271 3844
rect 5961 3776 6063 3810
rect 6097 3776 6135 3810
rect 6169 3776 6271 3810
rect 5961 3742 6271 3776
rect 5961 3708 6063 3742
rect 6097 3708 6135 3742
rect 6169 3708 6271 3742
rect 5961 3674 6271 3708
rect 5961 3640 6063 3674
rect 6097 3640 6135 3674
rect 6169 3640 6271 3674
rect 5961 3606 6271 3640
rect 5961 3572 6063 3606
rect 6097 3572 6135 3606
rect 6169 3572 6271 3606
rect 5961 3538 6271 3572
rect 5961 3504 6063 3538
rect 6097 3504 6135 3538
rect 6169 3504 6271 3538
rect 5961 3470 6271 3504
rect 5961 3436 6063 3470
rect 6097 3436 6135 3470
rect 6169 3436 6271 3470
rect 5961 3402 6271 3436
rect 5961 3368 6063 3402
rect 6097 3368 6135 3402
rect 6169 3368 6271 3402
rect 5961 3334 6271 3368
rect 5961 3300 6063 3334
rect 6097 3300 6135 3334
rect 6169 3300 6271 3334
rect 5961 3266 6271 3300
rect 5961 3232 6063 3266
rect 6097 3232 6135 3266
rect 6169 3232 6271 3266
rect 5961 3198 6271 3232
rect 5961 3164 6063 3198
rect 6097 3164 6135 3198
rect 6169 3164 6271 3198
rect 5961 3152 6271 3164
rect 6391 4082 6542 4152
rect 6682 4082 6833 4152
rect 6391 4048 6493 4082
rect 6527 4048 6542 4082
rect 6682 4048 6697 4082
rect 6731 4048 6833 4082
rect 6391 4014 6542 4048
rect 6682 4014 6833 4048
rect 6391 3980 6493 4014
rect 6527 3980 6542 4014
rect 6682 3980 6697 4014
rect 6731 3980 6833 4014
rect 6391 3946 6542 3980
rect 6682 3946 6833 3980
rect 6391 3912 6493 3946
rect 6527 3912 6542 3946
rect 6682 3912 6697 3946
rect 6731 3912 6833 3946
rect 6391 3878 6542 3912
rect 6682 3878 6833 3912
rect 6391 3844 6493 3878
rect 6527 3844 6542 3878
rect 6682 3844 6697 3878
rect 6731 3844 6833 3878
rect 6391 3810 6542 3844
rect 6682 3810 6833 3844
rect 6391 3776 6493 3810
rect 6527 3776 6542 3810
rect 6682 3776 6697 3810
rect 6731 3776 6833 3810
rect 6391 3742 6542 3776
rect 6682 3742 6833 3776
rect 6391 3708 6493 3742
rect 6527 3708 6542 3742
rect 6682 3708 6697 3742
rect 6731 3708 6833 3742
rect 6391 3674 6542 3708
rect 6682 3674 6833 3708
rect 6391 3640 6493 3674
rect 6527 3640 6542 3674
rect 6682 3640 6697 3674
rect 6731 3640 6833 3674
rect 6391 3606 6542 3640
rect 6682 3606 6833 3640
rect 6391 3572 6493 3606
rect 6527 3572 6542 3606
rect 6682 3572 6697 3606
rect 6731 3572 6833 3606
rect 6391 3538 6542 3572
rect 6682 3538 6833 3572
rect 6391 3504 6493 3538
rect 6527 3504 6542 3538
rect 6682 3504 6697 3538
rect 6731 3504 6833 3538
rect 6391 3470 6542 3504
rect 6682 3470 6833 3504
rect 6391 3436 6493 3470
rect 6527 3436 6542 3470
rect 6682 3436 6697 3470
rect 6731 3436 6833 3470
rect 6391 3402 6542 3436
rect 6682 3402 6833 3436
rect 6391 3368 6493 3402
rect 6527 3368 6542 3402
rect 6682 3368 6697 3402
rect 6731 3368 6833 3402
rect 6391 3334 6542 3368
rect 6682 3334 6833 3368
rect 6391 3300 6493 3334
rect 6527 3300 6542 3334
rect 6682 3300 6697 3334
rect 6731 3300 6833 3334
rect 6391 3266 6542 3300
rect 6682 3266 6833 3300
rect 6391 3232 6493 3266
rect 6527 3232 6542 3266
rect 6682 3232 6697 3266
rect 6731 3232 6833 3266
rect 6391 3198 6542 3232
rect 6682 3198 6833 3232
rect 6391 3164 6493 3198
rect 6527 3164 6542 3198
rect 6682 3164 6697 3198
rect 6731 3164 6833 3198
rect 6391 3152 6542 3164
rect 6682 3152 6833 3164
rect 6953 4082 7263 4152
rect 6953 4048 7055 4082
rect 7089 4048 7127 4082
rect 7161 4048 7263 4082
rect 6953 4014 7263 4048
rect 6953 3980 7055 4014
rect 7089 3980 7127 4014
rect 7161 3980 7263 4014
rect 6953 3946 7263 3980
rect 6953 3912 7055 3946
rect 7089 3912 7127 3946
rect 7161 3912 7263 3946
rect 6953 3878 7263 3912
rect 6953 3844 7055 3878
rect 7089 3844 7127 3878
rect 7161 3844 7263 3878
rect 6953 3810 7263 3844
rect 6953 3776 7055 3810
rect 7089 3776 7127 3810
rect 7161 3776 7263 3810
rect 6953 3742 7263 3776
rect 6953 3708 7055 3742
rect 7089 3708 7127 3742
rect 7161 3708 7263 3742
rect 6953 3674 7263 3708
rect 6953 3640 7055 3674
rect 7089 3640 7127 3674
rect 7161 3640 7263 3674
rect 6953 3606 7263 3640
rect 6953 3572 7055 3606
rect 7089 3572 7127 3606
rect 7161 3572 7263 3606
rect 6953 3538 7263 3572
rect 6953 3504 7055 3538
rect 7089 3504 7127 3538
rect 7161 3504 7263 3538
rect 6953 3470 7263 3504
rect 6953 3436 7055 3470
rect 7089 3436 7127 3470
rect 7161 3436 7263 3470
rect 6953 3402 7263 3436
rect 6953 3368 7055 3402
rect 7089 3368 7127 3402
rect 7161 3368 7263 3402
rect 6953 3334 7263 3368
rect 6953 3300 7055 3334
rect 7089 3300 7127 3334
rect 7161 3300 7263 3334
rect 6953 3266 7263 3300
rect 6953 3232 7055 3266
rect 7089 3232 7127 3266
rect 7161 3232 7263 3266
rect 6953 3198 7263 3232
rect 6953 3164 7055 3198
rect 7089 3164 7127 3198
rect 7161 3164 7263 3198
rect 6953 3152 7263 3164
rect 7383 4082 7534 4152
rect 7674 4082 7825 4152
rect 7383 4048 7485 4082
rect 7519 4048 7534 4082
rect 7674 4048 7689 4082
rect 7723 4048 7825 4082
rect 7383 4014 7534 4048
rect 7674 4014 7825 4048
rect 7383 3980 7485 4014
rect 7519 3980 7534 4014
rect 7674 3980 7689 4014
rect 7723 3980 7825 4014
rect 7383 3946 7534 3980
rect 7674 3946 7825 3980
rect 7383 3912 7485 3946
rect 7519 3912 7534 3946
rect 7674 3912 7689 3946
rect 7723 3912 7825 3946
rect 7383 3878 7534 3912
rect 7674 3878 7825 3912
rect 7383 3844 7485 3878
rect 7519 3844 7534 3878
rect 7674 3844 7689 3878
rect 7723 3844 7825 3878
rect 7383 3810 7534 3844
rect 7674 3810 7825 3844
rect 7383 3776 7485 3810
rect 7519 3776 7534 3810
rect 7674 3776 7689 3810
rect 7723 3776 7825 3810
rect 7383 3742 7534 3776
rect 7674 3742 7825 3776
rect 7383 3708 7485 3742
rect 7519 3708 7534 3742
rect 7674 3708 7689 3742
rect 7723 3708 7825 3742
rect 7383 3674 7534 3708
rect 7674 3674 7825 3708
rect 7383 3640 7485 3674
rect 7519 3640 7534 3674
rect 7674 3640 7689 3674
rect 7723 3640 7825 3674
rect 7383 3606 7534 3640
rect 7674 3606 7825 3640
rect 7383 3572 7485 3606
rect 7519 3572 7534 3606
rect 7674 3572 7689 3606
rect 7723 3572 7825 3606
rect 7383 3538 7534 3572
rect 7674 3538 7825 3572
rect 7383 3504 7485 3538
rect 7519 3504 7534 3538
rect 7674 3504 7689 3538
rect 7723 3504 7825 3538
rect 7383 3470 7534 3504
rect 7674 3470 7825 3504
rect 7383 3436 7485 3470
rect 7519 3436 7534 3470
rect 7674 3436 7689 3470
rect 7723 3436 7825 3470
rect 7383 3402 7534 3436
rect 7674 3402 7825 3436
rect 7383 3368 7485 3402
rect 7519 3368 7534 3402
rect 7674 3368 7689 3402
rect 7723 3368 7825 3402
rect 7383 3334 7534 3368
rect 7674 3334 7825 3368
rect 7383 3300 7485 3334
rect 7519 3300 7534 3334
rect 7674 3300 7689 3334
rect 7723 3300 7825 3334
rect 7383 3266 7534 3300
rect 7674 3266 7825 3300
rect 7383 3232 7485 3266
rect 7519 3232 7534 3266
rect 7674 3232 7689 3266
rect 7723 3232 7825 3266
rect 7383 3198 7534 3232
rect 7674 3198 7825 3232
rect 7383 3164 7485 3198
rect 7519 3164 7534 3198
rect 7674 3164 7689 3198
rect 7723 3164 7825 3198
rect 7383 3152 7534 3164
rect 7674 3152 7825 3164
rect 7945 4082 8255 4152
rect 7945 4048 8047 4082
rect 8081 4048 8119 4082
rect 8153 4048 8255 4082
rect 7945 4014 8255 4048
rect 7945 3980 8047 4014
rect 8081 3980 8119 4014
rect 8153 3980 8255 4014
rect 7945 3946 8255 3980
rect 7945 3912 8047 3946
rect 8081 3912 8119 3946
rect 8153 3912 8255 3946
rect 7945 3878 8255 3912
rect 7945 3844 8047 3878
rect 8081 3844 8119 3878
rect 8153 3844 8255 3878
rect 7945 3810 8255 3844
rect 7945 3776 8047 3810
rect 8081 3776 8119 3810
rect 8153 3776 8255 3810
rect 7945 3742 8255 3776
rect 7945 3708 8047 3742
rect 8081 3708 8119 3742
rect 8153 3708 8255 3742
rect 7945 3674 8255 3708
rect 7945 3640 8047 3674
rect 8081 3640 8119 3674
rect 8153 3640 8255 3674
rect 7945 3606 8255 3640
rect 7945 3572 8047 3606
rect 8081 3572 8119 3606
rect 8153 3572 8255 3606
rect 7945 3538 8255 3572
rect 7945 3504 8047 3538
rect 8081 3504 8119 3538
rect 8153 3504 8255 3538
rect 7945 3470 8255 3504
rect 7945 3436 8047 3470
rect 8081 3436 8119 3470
rect 8153 3436 8255 3470
rect 7945 3402 8255 3436
rect 7945 3368 8047 3402
rect 8081 3368 8119 3402
rect 8153 3368 8255 3402
rect 7945 3334 8255 3368
rect 7945 3300 8047 3334
rect 8081 3300 8119 3334
rect 8153 3300 8255 3334
rect 7945 3266 8255 3300
rect 7945 3232 8047 3266
rect 8081 3232 8119 3266
rect 8153 3232 8255 3266
rect 7945 3198 8255 3232
rect 7945 3164 8047 3198
rect 8081 3164 8119 3198
rect 8153 3164 8255 3198
rect 7945 3152 8255 3164
rect 8375 4082 8526 4152
rect 8666 4082 8817 4152
rect 8375 4048 8477 4082
rect 8511 4048 8526 4082
rect 8666 4048 8681 4082
rect 8715 4048 8817 4082
rect 8375 4014 8526 4048
rect 8666 4014 8817 4048
rect 8375 3980 8477 4014
rect 8511 3980 8526 4014
rect 8666 3980 8681 4014
rect 8715 3980 8817 4014
rect 8375 3946 8526 3980
rect 8666 3946 8817 3980
rect 8375 3912 8477 3946
rect 8511 3912 8526 3946
rect 8666 3912 8681 3946
rect 8715 3912 8817 3946
rect 8375 3878 8526 3912
rect 8666 3878 8817 3912
rect 8375 3844 8477 3878
rect 8511 3844 8526 3878
rect 8666 3844 8681 3878
rect 8715 3844 8817 3878
rect 8375 3810 8526 3844
rect 8666 3810 8817 3844
rect 8375 3776 8477 3810
rect 8511 3776 8526 3810
rect 8666 3776 8681 3810
rect 8715 3776 8817 3810
rect 8375 3742 8526 3776
rect 8666 3742 8817 3776
rect 8375 3708 8477 3742
rect 8511 3708 8526 3742
rect 8666 3708 8681 3742
rect 8715 3708 8817 3742
rect 8375 3674 8526 3708
rect 8666 3674 8817 3708
rect 8375 3640 8477 3674
rect 8511 3640 8526 3674
rect 8666 3640 8681 3674
rect 8715 3640 8817 3674
rect 8375 3606 8526 3640
rect 8666 3606 8817 3640
rect 8375 3572 8477 3606
rect 8511 3572 8526 3606
rect 8666 3572 8681 3606
rect 8715 3572 8817 3606
rect 8375 3538 8526 3572
rect 8666 3538 8817 3572
rect 8375 3504 8477 3538
rect 8511 3504 8526 3538
rect 8666 3504 8681 3538
rect 8715 3504 8817 3538
rect 8375 3470 8526 3504
rect 8666 3470 8817 3504
rect 8375 3436 8477 3470
rect 8511 3436 8526 3470
rect 8666 3436 8681 3470
rect 8715 3436 8817 3470
rect 8375 3402 8526 3436
rect 8666 3402 8817 3436
rect 8375 3368 8477 3402
rect 8511 3368 8526 3402
rect 8666 3368 8681 3402
rect 8715 3368 8817 3402
rect 8375 3334 8526 3368
rect 8666 3334 8817 3368
rect 8375 3300 8477 3334
rect 8511 3300 8526 3334
rect 8666 3300 8681 3334
rect 8715 3300 8817 3334
rect 8375 3266 8526 3300
rect 8666 3266 8817 3300
rect 8375 3232 8477 3266
rect 8511 3232 8526 3266
rect 8666 3232 8681 3266
rect 8715 3232 8817 3266
rect 8375 3198 8526 3232
rect 8666 3198 8817 3232
rect 8375 3164 8477 3198
rect 8511 3164 8526 3198
rect 8666 3164 8681 3198
rect 8715 3164 8817 3198
rect 8375 3152 8526 3164
rect 8666 3152 8817 3164
rect 8937 4082 9247 4152
rect 8937 4048 9039 4082
rect 9073 4048 9111 4082
rect 9145 4048 9247 4082
rect 8937 4014 9247 4048
rect 8937 3980 9039 4014
rect 9073 3980 9111 4014
rect 9145 3980 9247 4014
rect 8937 3946 9247 3980
rect 8937 3912 9039 3946
rect 9073 3912 9111 3946
rect 9145 3912 9247 3946
rect 8937 3878 9247 3912
rect 8937 3844 9039 3878
rect 9073 3844 9111 3878
rect 9145 3844 9247 3878
rect 8937 3810 9247 3844
rect 8937 3776 9039 3810
rect 9073 3776 9111 3810
rect 9145 3776 9247 3810
rect 8937 3742 9247 3776
rect 8937 3708 9039 3742
rect 9073 3708 9111 3742
rect 9145 3708 9247 3742
rect 8937 3674 9247 3708
rect 8937 3640 9039 3674
rect 9073 3640 9111 3674
rect 9145 3640 9247 3674
rect 8937 3606 9247 3640
rect 8937 3572 9039 3606
rect 9073 3572 9111 3606
rect 9145 3572 9247 3606
rect 8937 3538 9247 3572
rect 8937 3504 9039 3538
rect 9073 3504 9111 3538
rect 9145 3504 9247 3538
rect 8937 3470 9247 3504
rect 8937 3436 9039 3470
rect 9073 3436 9111 3470
rect 9145 3436 9247 3470
rect 8937 3402 9247 3436
rect 8937 3368 9039 3402
rect 9073 3368 9111 3402
rect 9145 3368 9247 3402
rect 8937 3334 9247 3368
rect 8937 3300 9039 3334
rect 9073 3300 9111 3334
rect 9145 3300 9247 3334
rect 8937 3266 9247 3300
rect 8937 3232 9039 3266
rect 9073 3232 9111 3266
rect 9145 3232 9247 3266
rect 8937 3198 9247 3232
rect 8937 3164 9039 3198
rect 9073 3164 9111 3198
rect 9145 3164 9247 3198
rect 8937 3152 9247 3164
rect 9367 4082 9518 4152
rect 9658 4082 9809 4152
rect 9367 4048 9469 4082
rect 9503 4048 9518 4082
rect 9658 4048 9673 4082
rect 9707 4048 9809 4082
rect 9367 4014 9518 4048
rect 9658 4014 9809 4048
rect 9367 3980 9469 4014
rect 9503 3980 9518 4014
rect 9658 3980 9673 4014
rect 9707 3980 9809 4014
rect 9367 3946 9518 3980
rect 9658 3946 9809 3980
rect 9367 3912 9469 3946
rect 9503 3912 9518 3946
rect 9658 3912 9673 3946
rect 9707 3912 9809 3946
rect 9367 3878 9518 3912
rect 9658 3878 9809 3912
rect 9367 3844 9469 3878
rect 9503 3844 9518 3878
rect 9658 3844 9673 3878
rect 9707 3844 9809 3878
rect 9367 3810 9518 3844
rect 9658 3810 9809 3844
rect 9367 3776 9469 3810
rect 9503 3776 9518 3810
rect 9658 3776 9673 3810
rect 9707 3776 9809 3810
rect 9367 3742 9518 3776
rect 9658 3742 9809 3776
rect 9367 3708 9469 3742
rect 9503 3708 9518 3742
rect 9658 3708 9673 3742
rect 9707 3708 9809 3742
rect 9367 3674 9518 3708
rect 9658 3674 9809 3708
rect 9367 3640 9469 3674
rect 9503 3640 9518 3674
rect 9658 3640 9673 3674
rect 9707 3640 9809 3674
rect 9367 3606 9518 3640
rect 9658 3606 9809 3640
rect 9367 3572 9469 3606
rect 9503 3572 9518 3606
rect 9658 3572 9673 3606
rect 9707 3572 9809 3606
rect 9367 3538 9518 3572
rect 9658 3538 9809 3572
rect 9367 3504 9469 3538
rect 9503 3504 9518 3538
rect 9658 3504 9673 3538
rect 9707 3504 9809 3538
rect 9367 3470 9518 3504
rect 9658 3470 9809 3504
rect 9367 3436 9469 3470
rect 9503 3436 9518 3470
rect 9658 3436 9673 3470
rect 9707 3436 9809 3470
rect 9367 3402 9518 3436
rect 9658 3402 9809 3436
rect 9367 3368 9469 3402
rect 9503 3368 9518 3402
rect 9658 3368 9673 3402
rect 9707 3368 9809 3402
rect 9367 3334 9518 3368
rect 9658 3334 9809 3368
rect 9367 3300 9469 3334
rect 9503 3300 9518 3334
rect 9658 3300 9673 3334
rect 9707 3300 9809 3334
rect 9367 3266 9518 3300
rect 9658 3266 9809 3300
rect 9367 3232 9469 3266
rect 9503 3232 9518 3266
rect 9658 3232 9673 3266
rect 9707 3232 9809 3266
rect 9367 3198 9518 3232
rect 9658 3198 9809 3232
rect 9367 3164 9469 3198
rect 9503 3164 9518 3198
rect 9658 3164 9673 3198
rect 9707 3164 9809 3198
rect 9367 3152 9518 3164
rect 9658 3152 9809 3164
rect 9929 4082 10239 4152
rect 9929 4048 10031 4082
rect 10065 4048 10103 4082
rect 10137 4048 10239 4082
rect 9929 4014 10239 4048
rect 9929 3980 10031 4014
rect 10065 3980 10103 4014
rect 10137 3980 10239 4014
rect 9929 3946 10239 3980
rect 9929 3912 10031 3946
rect 10065 3912 10103 3946
rect 10137 3912 10239 3946
rect 9929 3878 10239 3912
rect 9929 3844 10031 3878
rect 10065 3844 10103 3878
rect 10137 3844 10239 3878
rect 9929 3810 10239 3844
rect 9929 3776 10031 3810
rect 10065 3776 10103 3810
rect 10137 3776 10239 3810
rect 9929 3742 10239 3776
rect 9929 3708 10031 3742
rect 10065 3708 10103 3742
rect 10137 3708 10239 3742
rect 9929 3674 10239 3708
rect 9929 3640 10031 3674
rect 10065 3640 10103 3674
rect 10137 3640 10239 3674
rect 9929 3606 10239 3640
rect 9929 3572 10031 3606
rect 10065 3572 10103 3606
rect 10137 3572 10239 3606
rect 9929 3538 10239 3572
rect 9929 3504 10031 3538
rect 10065 3504 10103 3538
rect 10137 3504 10239 3538
rect 9929 3470 10239 3504
rect 9929 3436 10031 3470
rect 10065 3436 10103 3470
rect 10137 3436 10239 3470
rect 9929 3402 10239 3436
rect 9929 3368 10031 3402
rect 10065 3368 10103 3402
rect 10137 3368 10239 3402
rect 9929 3334 10239 3368
rect 9929 3300 10031 3334
rect 10065 3300 10103 3334
rect 10137 3300 10239 3334
rect 9929 3266 10239 3300
rect 9929 3232 10031 3266
rect 10065 3232 10103 3266
rect 10137 3232 10239 3266
rect 9929 3198 10239 3232
rect 9929 3164 10031 3198
rect 10065 3164 10103 3198
rect 10137 3164 10239 3198
rect 9929 3152 10239 3164
rect 10359 4082 10510 4152
rect 10650 4082 10801 4152
rect 10359 4048 10461 4082
rect 10495 4048 10510 4082
rect 10650 4048 10665 4082
rect 10699 4048 10801 4082
rect 10359 4014 10510 4048
rect 10650 4014 10801 4048
rect 10359 3980 10461 4014
rect 10495 3980 10510 4014
rect 10650 3980 10665 4014
rect 10699 3980 10801 4014
rect 10359 3946 10510 3980
rect 10650 3946 10801 3980
rect 10359 3912 10461 3946
rect 10495 3912 10510 3946
rect 10650 3912 10665 3946
rect 10699 3912 10801 3946
rect 10359 3878 10510 3912
rect 10650 3878 10801 3912
rect 10359 3844 10461 3878
rect 10495 3844 10510 3878
rect 10650 3844 10665 3878
rect 10699 3844 10801 3878
rect 10359 3810 10510 3844
rect 10650 3810 10801 3844
rect 10359 3776 10461 3810
rect 10495 3776 10510 3810
rect 10650 3776 10665 3810
rect 10699 3776 10801 3810
rect 10359 3742 10510 3776
rect 10650 3742 10801 3776
rect 10359 3708 10461 3742
rect 10495 3708 10510 3742
rect 10650 3708 10665 3742
rect 10699 3708 10801 3742
rect 10359 3674 10510 3708
rect 10650 3674 10801 3708
rect 10359 3640 10461 3674
rect 10495 3640 10510 3674
rect 10650 3640 10665 3674
rect 10699 3640 10801 3674
rect 10359 3606 10510 3640
rect 10650 3606 10801 3640
rect 10359 3572 10461 3606
rect 10495 3572 10510 3606
rect 10650 3572 10665 3606
rect 10699 3572 10801 3606
rect 10359 3538 10510 3572
rect 10650 3538 10801 3572
rect 10359 3504 10461 3538
rect 10495 3504 10510 3538
rect 10650 3504 10665 3538
rect 10699 3504 10801 3538
rect 10359 3470 10510 3504
rect 10650 3470 10801 3504
rect 10359 3436 10461 3470
rect 10495 3436 10510 3470
rect 10650 3436 10665 3470
rect 10699 3436 10801 3470
rect 10359 3402 10510 3436
rect 10650 3402 10801 3436
rect 10359 3368 10461 3402
rect 10495 3368 10510 3402
rect 10650 3368 10665 3402
rect 10699 3368 10801 3402
rect 10359 3334 10510 3368
rect 10650 3334 10801 3368
rect 10359 3300 10461 3334
rect 10495 3300 10510 3334
rect 10650 3300 10665 3334
rect 10699 3300 10801 3334
rect 10359 3266 10510 3300
rect 10650 3266 10801 3300
rect 10359 3232 10461 3266
rect 10495 3232 10510 3266
rect 10650 3232 10665 3266
rect 10699 3232 10801 3266
rect 10359 3198 10510 3232
rect 10650 3198 10801 3232
rect 10359 3164 10461 3198
rect 10495 3164 10510 3198
rect 10650 3164 10665 3198
rect 10699 3164 10801 3198
rect 10359 3152 10510 3164
rect 10650 3152 10801 3164
rect 10921 4082 11231 4152
rect 10921 4048 11023 4082
rect 11057 4048 11095 4082
rect 11129 4048 11231 4082
rect 10921 4014 11231 4048
rect 10921 3980 11023 4014
rect 11057 3980 11095 4014
rect 11129 3980 11231 4014
rect 10921 3946 11231 3980
rect 10921 3912 11023 3946
rect 11057 3912 11095 3946
rect 11129 3912 11231 3946
rect 10921 3878 11231 3912
rect 10921 3844 11023 3878
rect 11057 3844 11095 3878
rect 11129 3844 11231 3878
rect 10921 3810 11231 3844
rect 10921 3776 11023 3810
rect 11057 3776 11095 3810
rect 11129 3776 11231 3810
rect 10921 3742 11231 3776
rect 10921 3708 11023 3742
rect 11057 3708 11095 3742
rect 11129 3708 11231 3742
rect 10921 3674 11231 3708
rect 10921 3640 11023 3674
rect 11057 3640 11095 3674
rect 11129 3640 11231 3674
rect 10921 3606 11231 3640
rect 10921 3572 11023 3606
rect 11057 3572 11095 3606
rect 11129 3572 11231 3606
rect 10921 3538 11231 3572
rect 10921 3504 11023 3538
rect 11057 3504 11095 3538
rect 11129 3504 11231 3538
rect 10921 3470 11231 3504
rect 10921 3436 11023 3470
rect 11057 3436 11095 3470
rect 11129 3436 11231 3470
rect 10921 3402 11231 3436
rect 10921 3368 11023 3402
rect 11057 3368 11095 3402
rect 11129 3368 11231 3402
rect 10921 3334 11231 3368
rect 10921 3300 11023 3334
rect 11057 3300 11095 3334
rect 11129 3300 11231 3334
rect 10921 3266 11231 3300
rect 10921 3232 11023 3266
rect 11057 3232 11095 3266
rect 11129 3232 11231 3266
rect 10921 3198 11231 3232
rect 10921 3164 11023 3198
rect 11057 3164 11095 3198
rect 11129 3164 11231 3198
rect 10921 3152 11231 3164
rect 11351 4082 11502 4152
rect 11642 4082 11793 4152
rect 11351 4048 11453 4082
rect 11487 4048 11502 4082
rect 11642 4048 11657 4082
rect 11691 4048 11793 4082
rect 11351 4014 11502 4048
rect 11642 4014 11793 4048
rect 11351 3980 11453 4014
rect 11487 3980 11502 4014
rect 11642 3980 11657 4014
rect 11691 3980 11793 4014
rect 11351 3946 11502 3980
rect 11642 3946 11793 3980
rect 11351 3912 11453 3946
rect 11487 3912 11502 3946
rect 11642 3912 11657 3946
rect 11691 3912 11793 3946
rect 11351 3878 11502 3912
rect 11642 3878 11793 3912
rect 11351 3844 11453 3878
rect 11487 3844 11502 3878
rect 11642 3844 11657 3878
rect 11691 3844 11793 3878
rect 11351 3810 11502 3844
rect 11642 3810 11793 3844
rect 11351 3776 11453 3810
rect 11487 3776 11502 3810
rect 11642 3776 11657 3810
rect 11691 3776 11793 3810
rect 11351 3742 11502 3776
rect 11642 3742 11793 3776
rect 11351 3708 11453 3742
rect 11487 3708 11502 3742
rect 11642 3708 11657 3742
rect 11691 3708 11793 3742
rect 11351 3674 11502 3708
rect 11642 3674 11793 3708
rect 11351 3640 11453 3674
rect 11487 3640 11502 3674
rect 11642 3640 11657 3674
rect 11691 3640 11793 3674
rect 11351 3606 11502 3640
rect 11642 3606 11793 3640
rect 11351 3572 11453 3606
rect 11487 3572 11502 3606
rect 11642 3572 11657 3606
rect 11691 3572 11793 3606
rect 11351 3538 11502 3572
rect 11642 3538 11793 3572
rect 11351 3504 11453 3538
rect 11487 3504 11502 3538
rect 11642 3504 11657 3538
rect 11691 3504 11793 3538
rect 11351 3470 11502 3504
rect 11642 3470 11793 3504
rect 11351 3436 11453 3470
rect 11487 3436 11502 3470
rect 11642 3436 11657 3470
rect 11691 3436 11793 3470
rect 11351 3402 11502 3436
rect 11642 3402 11793 3436
rect 11351 3368 11453 3402
rect 11487 3368 11502 3402
rect 11642 3368 11657 3402
rect 11691 3368 11793 3402
rect 11351 3334 11502 3368
rect 11642 3334 11793 3368
rect 11351 3300 11453 3334
rect 11487 3300 11502 3334
rect 11642 3300 11657 3334
rect 11691 3300 11793 3334
rect 11351 3266 11502 3300
rect 11642 3266 11793 3300
rect 11351 3232 11453 3266
rect 11487 3232 11502 3266
rect 11642 3232 11657 3266
rect 11691 3232 11793 3266
rect 11351 3198 11502 3232
rect 11642 3198 11793 3232
rect 11351 3164 11453 3198
rect 11487 3164 11502 3198
rect 11642 3164 11657 3198
rect 11691 3164 11793 3198
rect 11351 3152 11502 3164
rect 11642 3152 11793 3164
rect 11913 4082 12223 4152
rect 11913 4048 12015 4082
rect 12049 4048 12087 4082
rect 12121 4048 12223 4082
rect 11913 4014 12223 4048
rect 11913 3980 12015 4014
rect 12049 3980 12087 4014
rect 12121 3980 12223 4014
rect 11913 3946 12223 3980
rect 11913 3912 12015 3946
rect 12049 3912 12087 3946
rect 12121 3912 12223 3946
rect 11913 3878 12223 3912
rect 11913 3844 12015 3878
rect 12049 3844 12087 3878
rect 12121 3844 12223 3878
rect 11913 3810 12223 3844
rect 11913 3776 12015 3810
rect 12049 3776 12087 3810
rect 12121 3776 12223 3810
rect 11913 3742 12223 3776
rect 11913 3708 12015 3742
rect 12049 3708 12087 3742
rect 12121 3708 12223 3742
rect 11913 3674 12223 3708
rect 11913 3640 12015 3674
rect 12049 3640 12087 3674
rect 12121 3640 12223 3674
rect 11913 3606 12223 3640
rect 11913 3572 12015 3606
rect 12049 3572 12087 3606
rect 12121 3572 12223 3606
rect 11913 3538 12223 3572
rect 11913 3504 12015 3538
rect 12049 3504 12087 3538
rect 12121 3504 12223 3538
rect 11913 3470 12223 3504
rect 11913 3436 12015 3470
rect 12049 3436 12087 3470
rect 12121 3436 12223 3470
rect 11913 3402 12223 3436
rect 11913 3368 12015 3402
rect 12049 3368 12087 3402
rect 12121 3368 12223 3402
rect 11913 3334 12223 3368
rect 11913 3300 12015 3334
rect 12049 3300 12087 3334
rect 12121 3300 12223 3334
rect 11913 3266 12223 3300
rect 11913 3232 12015 3266
rect 12049 3232 12087 3266
rect 12121 3232 12223 3266
rect 11913 3198 12223 3232
rect 11913 3164 12015 3198
rect 12049 3164 12087 3198
rect 12121 3164 12223 3198
rect 11913 3152 12223 3164
rect 12343 4082 12494 4152
rect 12634 4082 12785 4152
rect 12343 4048 12445 4082
rect 12479 4048 12494 4082
rect 12634 4048 12649 4082
rect 12683 4048 12785 4082
rect 12343 4014 12494 4048
rect 12634 4014 12785 4048
rect 12343 3980 12445 4014
rect 12479 3980 12494 4014
rect 12634 3980 12649 4014
rect 12683 3980 12785 4014
rect 12343 3946 12494 3980
rect 12634 3946 12785 3980
rect 12343 3912 12445 3946
rect 12479 3912 12494 3946
rect 12634 3912 12649 3946
rect 12683 3912 12785 3946
rect 12343 3878 12494 3912
rect 12634 3878 12785 3912
rect 12343 3844 12445 3878
rect 12479 3844 12494 3878
rect 12634 3844 12649 3878
rect 12683 3844 12785 3878
rect 12343 3810 12494 3844
rect 12634 3810 12785 3844
rect 12343 3776 12445 3810
rect 12479 3776 12494 3810
rect 12634 3776 12649 3810
rect 12683 3776 12785 3810
rect 12343 3742 12494 3776
rect 12634 3742 12785 3776
rect 12343 3708 12445 3742
rect 12479 3708 12494 3742
rect 12634 3708 12649 3742
rect 12683 3708 12785 3742
rect 12343 3674 12494 3708
rect 12634 3674 12785 3708
rect 12343 3640 12445 3674
rect 12479 3640 12494 3674
rect 12634 3640 12649 3674
rect 12683 3640 12785 3674
rect 12343 3606 12494 3640
rect 12634 3606 12785 3640
rect 12343 3572 12445 3606
rect 12479 3572 12494 3606
rect 12634 3572 12649 3606
rect 12683 3572 12785 3606
rect 12343 3538 12494 3572
rect 12634 3538 12785 3572
rect 12343 3504 12445 3538
rect 12479 3504 12494 3538
rect 12634 3504 12649 3538
rect 12683 3504 12785 3538
rect 12343 3470 12494 3504
rect 12634 3470 12785 3504
rect 12343 3436 12445 3470
rect 12479 3436 12494 3470
rect 12634 3436 12649 3470
rect 12683 3436 12785 3470
rect 12343 3402 12494 3436
rect 12634 3402 12785 3436
rect 12343 3368 12445 3402
rect 12479 3368 12494 3402
rect 12634 3368 12649 3402
rect 12683 3368 12785 3402
rect 12343 3334 12494 3368
rect 12634 3334 12785 3368
rect 12343 3300 12445 3334
rect 12479 3300 12494 3334
rect 12634 3300 12649 3334
rect 12683 3300 12785 3334
rect 12343 3266 12494 3300
rect 12634 3266 12785 3300
rect 12343 3232 12445 3266
rect 12479 3232 12494 3266
rect 12634 3232 12649 3266
rect 12683 3232 12785 3266
rect 12343 3198 12494 3232
rect 12634 3198 12785 3232
rect 12343 3164 12445 3198
rect 12479 3164 12494 3198
rect 12634 3164 12649 3198
rect 12683 3164 12785 3198
rect 12343 3152 12494 3164
rect 12634 3152 12785 3164
rect 12905 4082 13215 4152
rect 12905 4048 13007 4082
rect 13041 4048 13079 4082
rect 13113 4048 13215 4082
rect 12905 4014 13215 4048
rect 12905 3980 13007 4014
rect 13041 3980 13079 4014
rect 13113 3980 13215 4014
rect 12905 3946 13215 3980
rect 12905 3912 13007 3946
rect 13041 3912 13079 3946
rect 13113 3912 13215 3946
rect 12905 3878 13215 3912
rect 12905 3844 13007 3878
rect 13041 3844 13079 3878
rect 13113 3844 13215 3878
rect 12905 3810 13215 3844
rect 12905 3776 13007 3810
rect 13041 3776 13079 3810
rect 13113 3776 13215 3810
rect 12905 3742 13215 3776
rect 12905 3708 13007 3742
rect 13041 3708 13079 3742
rect 13113 3708 13215 3742
rect 12905 3674 13215 3708
rect 12905 3640 13007 3674
rect 13041 3640 13079 3674
rect 13113 3640 13215 3674
rect 12905 3606 13215 3640
rect 12905 3572 13007 3606
rect 13041 3572 13079 3606
rect 13113 3572 13215 3606
rect 12905 3538 13215 3572
rect 12905 3504 13007 3538
rect 13041 3504 13079 3538
rect 13113 3504 13215 3538
rect 12905 3470 13215 3504
rect 12905 3436 13007 3470
rect 13041 3436 13079 3470
rect 13113 3436 13215 3470
rect 12905 3402 13215 3436
rect 12905 3368 13007 3402
rect 13041 3368 13079 3402
rect 13113 3368 13215 3402
rect 12905 3334 13215 3368
rect 12905 3300 13007 3334
rect 13041 3300 13079 3334
rect 13113 3300 13215 3334
rect 12905 3266 13215 3300
rect 12905 3232 13007 3266
rect 13041 3232 13079 3266
rect 13113 3232 13215 3266
rect 12905 3198 13215 3232
rect 12905 3164 13007 3198
rect 13041 3164 13079 3198
rect 13113 3164 13215 3198
rect 12905 3152 13215 3164
rect 13335 4082 13486 4152
rect 13626 4082 13777 4152
rect 13335 4048 13437 4082
rect 13471 4048 13486 4082
rect 13626 4048 13641 4082
rect 13675 4048 13777 4082
rect 13335 4014 13486 4048
rect 13626 4014 13777 4048
rect 13335 3980 13437 4014
rect 13471 3980 13486 4014
rect 13626 3980 13641 4014
rect 13675 3980 13777 4014
rect 13335 3946 13486 3980
rect 13626 3946 13777 3980
rect 13335 3912 13437 3946
rect 13471 3912 13486 3946
rect 13626 3912 13641 3946
rect 13675 3912 13777 3946
rect 13335 3878 13486 3912
rect 13626 3878 13777 3912
rect 13335 3844 13437 3878
rect 13471 3844 13486 3878
rect 13626 3844 13641 3878
rect 13675 3844 13777 3878
rect 13335 3810 13486 3844
rect 13626 3810 13777 3844
rect 13335 3776 13437 3810
rect 13471 3776 13486 3810
rect 13626 3776 13641 3810
rect 13675 3776 13777 3810
rect 13335 3742 13486 3776
rect 13626 3742 13777 3776
rect 13335 3708 13437 3742
rect 13471 3708 13486 3742
rect 13626 3708 13641 3742
rect 13675 3708 13777 3742
rect 13335 3674 13486 3708
rect 13626 3674 13777 3708
rect 13335 3640 13437 3674
rect 13471 3640 13486 3674
rect 13626 3640 13641 3674
rect 13675 3640 13777 3674
rect 13335 3606 13486 3640
rect 13626 3606 13777 3640
rect 13335 3572 13437 3606
rect 13471 3572 13486 3606
rect 13626 3572 13641 3606
rect 13675 3572 13777 3606
rect 13335 3538 13486 3572
rect 13626 3538 13777 3572
rect 13335 3504 13437 3538
rect 13471 3504 13486 3538
rect 13626 3504 13641 3538
rect 13675 3504 13777 3538
rect 13335 3470 13486 3504
rect 13626 3470 13777 3504
rect 13335 3436 13437 3470
rect 13471 3436 13486 3470
rect 13626 3436 13641 3470
rect 13675 3436 13777 3470
rect 13335 3402 13486 3436
rect 13626 3402 13777 3436
rect 13335 3368 13437 3402
rect 13471 3368 13486 3402
rect 13626 3368 13641 3402
rect 13675 3368 13777 3402
rect 13335 3334 13486 3368
rect 13626 3334 13777 3368
rect 13335 3300 13437 3334
rect 13471 3300 13486 3334
rect 13626 3300 13641 3334
rect 13675 3300 13777 3334
rect 13335 3266 13486 3300
rect 13626 3266 13777 3300
rect 13335 3232 13437 3266
rect 13471 3232 13486 3266
rect 13626 3232 13641 3266
rect 13675 3232 13777 3266
rect 13335 3198 13486 3232
rect 13626 3198 13777 3232
rect 13335 3164 13437 3198
rect 13471 3164 13486 3198
rect 13626 3164 13641 3198
rect 13675 3164 13777 3198
rect 13335 3152 13486 3164
rect 13626 3152 13777 3164
rect 13897 4082 14135 4152
rect 13897 4048 13999 4082
rect 14033 4048 14135 4082
rect 13897 4014 14135 4048
rect 13897 3980 13999 4014
rect 14033 3980 14135 4014
rect 13897 3946 14135 3980
rect 13897 3912 13999 3946
rect 14033 3912 14135 3946
rect 13897 3878 14135 3912
rect 13897 3844 13999 3878
rect 14033 3844 14135 3878
rect 13897 3810 14135 3844
rect 13897 3776 13999 3810
rect 14033 3776 14135 3810
rect 13897 3742 14135 3776
rect 13897 3708 13999 3742
rect 14033 3708 14135 3742
rect 13897 3674 14135 3708
rect 13897 3640 13999 3674
rect 14033 3640 14135 3674
rect 13897 3606 14135 3640
rect 13897 3572 13999 3606
rect 14033 3572 14135 3606
rect 13897 3538 14135 3572
rect 13897 3504 13999 3538
rect 14033 3504 14135 3538
rect 13897 3470 14135 3504
rect 13897 3436 13999 3470
rect 14033 3436 14135 3470
rect 13897 3402 14135 3436
rect 13897 3368 13999 3402
rect 14033 3368 14135 3402
rect 13897 3334 14135 3368
rect 13897 3300 13999 3334
rect 14033 3300 14135 3334
rect 13897 3266 14135 3300
rect 13897 3232 13999 3266
rect 14033 3232 14135 3266
rect 13897 3198 14135 3232
rect 13897 3164 13999 3198
rect 14033 3164 14135 3198
rect 13897 3152 14135 3164
rect 14255 4082 14427 4152
rect 14255 4048 14356 4082
rect 14390 4048 14427 4082
rect 14255 4014 14427 4048
rect 14255 3980 14356 4014
rect 14390 3980 14427 4014
rect 14255 3946 14427 3980
rect 14255 3912 14356 3946
rect 14390 3912 14427 3946
rect 14255 3878 14427 3912
rect 14255 3844 14356 3878
rect 14390 3844 14427 3878
rect 14255 3810 14427 3844
rect 14255 3776 14356 3810
rect 14390 3776 14427 3810
rect 14255 3742 14427 3776
rect 14255 3708 14356 3742
rect 14390 3708 14427 3742
rect 14255 3674 14427 3708
rect 14255 3640 14356 3674
rect 14390 3640 14427 3674
rect 14255 3606 14427 3640
rect 14255 3572 14356 3606
rect 14390 3572 14427 3606
rect 14255 3538 14427 3572
rect 14255 3504 14356 3538
rect 14390 3504 14427 3538
rect 14255 3470 14427 3504
rect 14255 3436 14356 3470
rect 14390 3436 14427 3470
rect 14255 3402 14427 3436
rect 14255 3368 14356 3402
rect 14390 3368 14427 3402
rect 14255 3334 14427 3368
rect 14255 3300 14356 3334
rect 14390 3300 14427 3334
rect 14255 3266 14427 3300
rect 14255 3232 14356 3266
rect 14390 3232 14427 3266
rect 14255 3198 14427 3232
rect 14255 3164 14356 3198
rect 14390 3164 14427 3198
rect 14255 3152 14427 3164
rect 708 2482 881 2552
rect 708 2448 745 2482
rect 779 2448 881 2482
rect 708 2414 881 2448
rect 708 2380 745 2414
rect 779 2380 881 2414
rect 708 2346 881 2380
rect 708 2312 745 2346
rect 779 2312 881 2346
rect 708 2278 881 2312
rect 708 2244 745 2278
rect 779 2244 881 2278
rect 708 2210 881 2244
rect 708 2176 745 2210
rect 779 2176 881 2210
rect 708 2142 881 2176
rect 708 2108 745 2142
rect 779 2108 881 2142
rect 708 2074 881 2108
rect 708 2040 745 2074
rect 779 2040 881 2074
rect 708 2006 881 2040
rect 708 1972 745 2006
rect 779 1972 881 2006
rect 708 1938 881 1972
rect 708 1904 745 1938
rect 779 1904 881 1938
rect 708 1870 881 1904
rect 708 1836 745 1870
rect 779 1836 881 1870
rect 708 1802 881 1836
rect 708 1768 745 1802
rect 779 1768 881 1802
rect 708 1734 881 1768
rect 708 1700 745 1734
rect 779 1700 881 1734
rect 708 1666 881 1700
rect 708 1632 745 1666
rect 779 1632 881 1666
rect 708 1598 881 1632
rect 708 1564 745 1598
rect 779 1564 881 1598
rect 708 1552 881 1564
rect 1001 2482 1311 2552
rect 1001 2448 1103 2482
rect 1137 2448 1175 2482
rect 1209 2448 1311 2482
rect 1001 2414 1311 2448
rect 1001 2380 1103 2414
rect 1137 2380 1175 2414
rect 1209 2380 1311 2414
rect 1001 2346 1311 2380
rect 1001 2312 1103 2346
rect 1137 2312 1175 2346
rect 1209 2312 1311 2346
rect 1001 2278 1311 2312
rect 1001 2244 1103 2278
rect 1137 2244 1175 2278
rect 1209 2244 1311 2278
rect 1001 2210 1311 2244
rect 1001 2176 1103 2210
rect 1137 2176 1175 2210
rect 1209 2176 1311 2210
rect 1001 2142 1311 2176
rect 1001 2108 1103 2142
rect 1137 2108 1175 2142
rect 1209 2108 1311 2142
rect 1001 2074 1311 2108
rect 1001 2040 1103 2074
rect 1137 2040 1175 2074
rect 1209 2040 1311 2074
rect 1001 2006 1311 2040
rect 1001 1972 1103 2006
rect 1137 1972 1175 2006
rect 1209 1972 1311 2006
rect 1001 1938 1311 1972
rect 1001 1904 1103 1938
rect 1137 1904 1175 1938
rect 1209 1904 1311 1938
rect 1001 1870 1311 1904
rect 1001 1836 1103 1870
rect 1137 1836 1175 1870
rect 1209 1836 1311 1870
rect 1001 1802 1311 1836
rect 1001 1768 1103 1802
rect 1137 1768 1175 1802
rect 1209 1768 1311 1802
rect 1001 1734 1311 1768
rect 1001 1700 1103 1734
rect 1137 1700 1175 1734
rect 1209 1700 1311 1734
rect 1001 1666 1311 1700
rect 1001 1632 1103 1666
rect 1137 1632 1175 1666
rect 1209 1632 1311 1666
rect 1001 1598 1311 1632
rect 1001 1564 1103 1598
rect 1137 1564 1175 1598
rect 1209 1564 1311 1598
rect 1001 1552 1311 1564
rect 1431 2540 1582 2552
rect 1722 2540 1873 2552
rect 1431 2506 1533 2540
rect 1567 2506 1582 2540
rect 1722 2506 1737 2540
rect 1771 2506 1873 2540
rect 1431 2472 1582 2506
rect 1722 2472 1873 2506
rect 1431 2438 1533 2472
rect 1567 2438 1582 2472
rect 1722 2438 1737 2472
rect 1771 2438 1873 2472
rect 1431 2404 1582 2438
rect 1722 2404 1873 2438
rect 1431 2370 1533 2404
rect 1567 2370 1582 2404
rect 1722 2370 1737 2404
rect 1771 2370 1873 2404
rect 1431 2336 1582 2370
rect 1722 2336 1873 2370
rect 1431 2302 1533 2336
rect 1567 2302 1582 2336
rect 1722 2302 1737 2336
rect 1771 2302 1873 2336
rect 1431 2268 1582 2302
rect 1722 2268 1873 2302
rect 1431 2234 1533 2268
rect 1567 2234 1582 2268
rect 1722 2234 1737 2268
rect 1771 2234 1873 2268
rect 1431 2200 1582 2234
rect 1722 2200 1873 2234
rect 1431 2166 1533 2200
rect 1567 2166 1582 2200
rect 1722 2166 1737 2200
rect 1771 2166 1873 2200
rect 1431 2132 1582 2166
rect 1722 2132 1873 2166
rect 1431 2098 1533 2132
rect 1567 2098 1582 2132
rect 1722 2098 1737 2132
rect 1771 2098 1873 2132
rect 1431 2064 1582 2098
rect 1722 2064 1873 2098
rect 1431 2030 1533 2064
rect 1567 2030 1582 2064
rect 1722 2030 1737 2064
rect 1771 2030 1873 2064
rect 1431 1996 1582 2030
rect 1722 1996 1873 2030
rect 1431 1962 1533 1996
rect 1567 1962 1582 1996
rect 1722 1962 1737 1996
rect 1771 1962 1873 1996
rect 1431 1928 1582 1962
rect 1722 1928 1873 1962
rect 1431 1894 1533 1928
rect 1567 1894 1582 1928
rect 1722 1894 1737 1928
rect 1771 1894 1873 1928
rect 1431 1860 1582 1894
rect 1722 1860 1873 1894
rect 1431 1826 1533 1860
rect 1567 1826 1582 1860
rect 1722 1826 1737 1860
rect 1771 1826 1873 1860
rect 1431 1792 1582 1826
rect 1722 1792 1873 1826
rect 1431 1758 1533 1792
rect 1567 1758 1582 1792
rect 1722 1758 1737 1792
rect 1771 1758 1873 1792
rect 1431 1724 1582 1758
rect 1722 1724 1873 1758
rect 1431 1690 1533 1724
rect 1567 1690 1582 1724
rect 1722 1690 1737 1724
rect 1771 1690 1873 1724
rect 1431 1656 1582 1690
rect 1722 1656 1873 1690
rect 1431 1622 1533 1656
rect 1567 1622 1582 1656
rect 1722 1622 1737 1656
rect 1771 1622 1873 1656
rect 1431 1552 1582 1622
rect 1722 1552 1873 1622
rect 1993 2482 2303 2552
rect 1993 2448 2095 2482
rect 2129 2448 2167 2482
rect 2201 2448 2303 2482
rect 1993 2414 2303 2448
rect 1993 2380 2095 2414
rect 2129 2380 2167 2414
rect 2201 2380 2303 2414
rect 1993 2346 2303 2380
rect 1993 2312 2095 2346
rect 2129 2312 2167 2346
rect 2201 2312 2303 2346
rect 1993 2278 2303 2312
rect 1993 2244 2095 2278
rect 2129 2244 2167 2278
rect 2201 2244 2303 2278
rect 1993 2210 2303 2244
rect 1993 2176 2095 2210
rect 2129 2176 2167 2210
rect 2201 2176 2303 2210
rect 1993 2142 2303 2176
rect 1993 2108 2095 2142
rect 2129 2108 2167 2142
rect 2201 2108 2303 2142
rect 1993 2074 2303 2108
rect 1993 2040 2095 2074
rect 2129 2040 2167 2074
rect 2201 2040 2303 2074
rect 1993 2006 2303 2040
rect 1993 1972 2095 2006
rect 2129 1972 2167 2006
rect 2201 1972 2303 2006
rect 1993 1938 2303 1972
rect 1993 1904 2095 1938
rect 2129 1904 2167 1938
rect 2201 1904 2303 1938
rect 1993 1870 2303 1904
rect 1993 1836 2095 1870
rect 2129 1836 2167 1870
rect 2201 1836 2303 1870
rect 1993 1802 2303 1836
rect 1993 1768 2095 1802
rect 2129 1768 2167 1802
rect 2201 1768 2303 1802
rect 1993 1734 2303 1768
rect 1993 1700 2095 1734
rect 2129 1700 2167 1734
rect 2201 1700 2303 1734
rect 1993 1666 2303 1700
rect 1993 1632 2095 1666
rect 2129 1632 2167 1666
rect 2201 1632 2303 1666
rect 1993 1598 2303 1632
rect 1993 1564 2095 1598
rect 2129 1564 2167 1598
rect 2201 1564 2303 1598
rect 1993 1552 2303 1564
rect 2423 2540 2574 2552
rect 2714 2540 2865 2552
rect 2423 2506 2525 2540
rect 2559 2506 2574 2540
rect 2714 2506 2729 2540
rect 2763 2506 2865 2540
rect 2423 2472 2574 2506
rect 2714 2472 2865 2506
rect 2423 2438 2525 2472
rect 2559 2438 2574 2472
rect 2714 2438 2729 2472
rect 2763 2438 2865 2472
rect 2423 2404 2574 2438
rect 2714 2404 2865 2438
rect 2423 2370 2525 2404
rect 2559 2370 2574 2404
rect 2714 2370 2729 2404
rect 2763 2370 2865 2404
rect 2423 2336 2574 2370
rect 2714 2336 2865 2370
rect 2423 2302 2525 2336
rect 2559 2302 2574 2336
rect 2714 2302 2729 2336
rect 2763 2302 2865 2336
rect 2423 2268 2574 2302
rect 2714 2268 2865 2302
rect 2423 2234 2525 2268
rect 2559 2234 2574 2268
rect 2714 2234 2729 2268
rect 2763 2234 2865 2268
rect 2423 2200 2574 2234
rect 2714 2200 2865 2234
rect 2423 2166 2525 2200
rect 2559 2166 2574 2200
rect 2714 2166 2729 2200
rect 2763 2166 2865 2200
rect 2423 2132 2574 2166
rect 2714 2132 2865 2166
rect 2423 2098 2525 2132
rect 2559 2098 2574 2132
rect 2714 2098 2729 2132
rect 2763 2098 2865 2132
rect 2423 2064 2574 2098
rect 2714 2064 2865 2098
rect 2423 2030 2525 2064
rect 2559 2030 2574 2064
rect 2714 2030 2729 2064
rect 2763 2030 2865 2064
rect 2423 1996 2574 2030
rect 2714 1996 2865 2030
rect 2423 1962 2525 1996
rect 2559 1962 2574 1996
rect 2714 1962 2729 1996
rect 2763 1962 2865 1996
rect 2423 1928 2574 1962
rect 2714 1928 2865 1962
rect 2423 1894 2525 1928
rect 2559 1894 2574 1928
rect 2714 1894 2729 1928
rect 2763 1894 2865 1928
rect 2423 1860 2574 1894
rect 2714 1860 2865 1894
rect 2423 1826 2525 1860
rect 2559 1826 2574 1860
rect 2714 1826 2729 1860
rect 2763 1826 2865 1860
rect 2423 1792 2574 1826
rect 2714 1792 2865 1826
rect 2423 1758 2525 1792
rect 2559 1758 2574 1792
rect 2714 1758 2729 1792
rect 2763 1758 2865 1792
rect 2423 1724 2574 1758
rect 2714 1724 2865 1758
rect 2423 1690 2525 1724
rect 2559 1690 2574 1724
rect 2714 1690 2729 1724
rect 2763 1690 2865 1724
rect 2423 1656 2574 1690
rect 2714 1656 2865 1690
rect 2423 1622 2525 1656
rect 2559 1622 2574 1656
rect 2714 1622 2729 1656
rect 2763 1622 2865 1656
rect 2423 1552 2574 1622
rect 2714 1552 2865 1622
rect 2985 2482 3295 2552
rect 2985 2448 3087 2482
rect 3121 2448 3159 2482
rect 3193 2448 3295 2482
rect 2985 2414 3295 2448
rect 2985 2380 3087 2414
rect 3121 2380 3159 2414
rect 3193 2380 3295 2414
rect 2985 2346 3295 2380
rect 2985 2312 3087 2346
rect 3121 2312 3159 2346
rect 3193 2312 3295 2346
rect 2985 2278 3295 2312
rect 2985 2244 3087 2278
rect 3121 2244 3159 2278
rect 3193 2244 3295 2278
rect 2985 2210 3295 2244
rect 2985 2176 3087 2210
rect 3121 2176 3159 2210
rect 3193 2176 3295 2210
rect 2985 2142 3295 2176
rect 2985 2108 3087 2142
rect 3121 2108 3159 2142
rect 3193 2108 3295 2142
rect 2985 2074 3295 2108
rect 2985 2040 3087 2074
rect 3121 2040 3159 2074
rect 3193 2040 3295 2074
rect 2985 2006 3295 2040
rect 2985 1972 3087 2006
rect 3121 1972 3159 2006
rect 3193 1972 3295 2006
rect 2985 1938 3295 1972
rect 2985 1904 3087 1938
rect 3121 1904 3159 1938
rect 3193 1904 3295 1938
rect 2985 1870 3295 1904
rect 2985 1836 3087 1870
rect 3121 1836 3159 1870
rect 3193 1836 3295 1870
rect 2985 1802 3295 1836
rect 2985 1768 3087 1802
rect 3121 1768 3159 1802
rect 3193 1768 3295 1802
rect 2985 1734 3295 1768
rect 2985 1700 3087 1734
rect 3121 1700 3159 1734
rect 3193 1700 3295 1734
rect 2985 1666 3295 1700
rect 2985 1632 3087 1666
rect 3121 1632 3159 1666
rect 3193 1632 3295 1666
rect 2985 1598 3295 1632
rect 2985 1564 3087 1598
rect 3121 1564 3159 1598
rect 3193 1564 3295 1598
rect 2985 1552 3295 1564
rect 3415 2540 3566 2552
rect 3706 2540 3857 2552
rect 3415 2506 3517 2540
rect 3551 2506 3566 2540
rect 3706 2506 3721 2540
rect 3755 2506 3857 2540
rect 3415 2472 3566 2506
rect 3706 2472 3857 2506
rect 3415 2438 3517 2472
rect 3551 2438 3566 2472
rect 3706 2438 3721 2472
rect 3755 2438 3857 2472
rect 3415 2404 3566 2438
rect 3706 2404 3857 2438
rect 3415 2370 3517 2404
rect 3551 2370 3566 2404
rect 3706 2370 3721 2404
rect 3755 2370 3857 2404
rect 3415 2336 3566 2370
rect 3706 2336 3857 2370
rect 3415 2302 3517 2336
rect 3551 2302 3566 2336
rect 3706 2302 3721 2336
rect 3755 2302 3857 2336
rect 3415 2268 3566 2302
rect 3706 2268 3857 2302
rect 3415 2234 3517 2268
rect 3551 2234 3566 2268
rect 3706 2234 3721 2268
rect 3755 2234 3857 2268
rect 3415 2200 3566 2234
rect 3706 2200 3857 2234
rect 3415 2166 3517 2200
rect 3551 2166 3566 2200
rect 3706 2166 3721 2200
rect 3755 2166 3857 2200
rect 3415 2132 3566 2166
rect 3706 2132 3857 2166
rect 3415 2098 3517 2132
rect 3551 2098 3566 2132
rect 3706 2098 3721 2132
rect 3755 2098 3857 2132
rect 3415 2064 3566 2098
rect 3706 2064 3857 2098
rect 3415 2030 3517 2064
rect 3551 2030 3566 2064
rect 3706 2030 3721 2064
rect 3755 2030 3857 2064
rect 3415 1996 3566 2030
rect 3706 1996 3857 2030
rect 3415 1962 3517 1996
rect 3551 1962 3566 1996
rect 3706 1962 3721 1996
rect 3755 1962 3857 1996
rect 3415 1928 3566 1962
rect 3706 1928 3857 1962
rect 3415 1894 3517 1928
rect 3551 1894 3566 1928
rect 3706 1894 3721 1928
rect 3755 1894 3857 1928
rect 3415 1860 3566 1894
rect 3706 1860 3857 1894
rect 3415 1826 3517 1860
rect 3551 1826 3566 1860
rect 3706 1826 3721 1860
rect 3755 1826 3857 1860
rect 3415 1792 3566 1826
rect 3706 1792 3857 1826
rect 3415 1758 3517 1792
rect 3551 1758 3566 1792
rect 3706 1758 3721 1792
rect 3755 1758 3857 1792
rect 3415 1724 3566 1758
rect 3706 1724 3857 1758
rect 3415 1690 3517 1724
rect 3551 1690 3566 1724
rect 3706 1690 3721 1724
rect 3755 1690 3857 1724
rect 3415 1656 3566 1690
rect 3706 1656 3857 1690
rect 3415 1622 3517 1656
rect 3551 1622 3566 1656
rect 3706 1622 3721 1656
rect 3755 1622 3857 1656
rect 3415 1552 3566 1622
rect 3706 1552 3857 1622
rect 3977 2482 4287 2552
rect 3977 2448 4079 2482
rect 4113 2448 4151 2482
rect 4185 2448 4287 2482
rect 3977 2414 4287 2448
rect 3977 2380 4079 2414
rect 4113 2380 4151 2414
rect 4185 2380 4287 2414
rect 3977 2346 4287 2380
rect 3977 2312 4079 2346
rect 4113 2312 4151 2346
rect 4185 2312 4287 2346
rect 3977 2278 4287 2312
rect 3977 2244 4079 2278
rect 4113 2244 4151 2278
rect 4185 2244 4287 2278
rect 3977 2210 4287 2244
rect 3977 2176 4079 2210
rect 4113 2176 4151 2210
rect 4185 2176 4287 2210
rect 3977 2142 4287 2176
rect 3977 2108 4079 2142
rect 4113 2108 4151 2142
rect 4185 2108 4287 2142
rect 3977 2074 4287 2108
rect 3977 2040 4079 2074
rect 4113 2040 4151 2074
rect 4185 2040 4287 2074
rect 3977 2006 4287 2040
rect 3977 1972 4079 2006
rect 4113 1972 4151 2006
rect 4185 1972 4287 2006
rect 3977 1938 4287 1972
rect 3977 1904 4079 1938
rect 4113 1904 4151 1938
rect 4185 1904 4287 1938
rect 3977 1870 4287 1904
rect 3977 1836 4079 1870
rect 4113 1836 4151 1870
rect 4185 1836 4287 1870
rect 3977 1802 4287 1836
rect 3977 1768 4079 1802
rect 4113 1768 4151 1802
rect 4185 1768 4287 1802
rect 3977 1734 4287 1768
rect 3977 1700 4079 1734
rect 4113 1700 4151 1734
rect 4185 1700 4287 1734
rect 3977 1666 4287 1700
rect 3977 1632 4079 1666
rect 4113 1632 4151 1666
rect 4185 1632 4287 1666
rect 3977 1598 4287 1632
rect 3977 1564 4079 1598
rect 4113 1564 4151 1598
rect 4185 1564 4287 1598
rect 3977 1552 4287 1564
rect 4407 2540 4558 2552
rect 4698 2540 4849 2552
rect 4407 2506 4509 2540
rect 4543 2506 4558 2540
rect 4698 2506 4713 2540
rect 4747 2506 4849 2540
rect 4407 2472 4558 2506
rect 4698 2472 4849 2506
rect 4407 2438 4509 2472
rect 4543 2438 4558 2472
rect 4698 2438 4713 2472
rect 4747 2438 4849 2472
rect 4407 2404 4558 2438
rect 4698 2404 4849 2438
rect 4407 2370 4509 2404
rect 4543 2370 4558 2404
rect 4698 2370 4713 2404
rect 4747 2370 4849 2404
rect 4407 2336 4558 2370
rect 4698 2336 4849 2370
rect 4407 2302 4509 2336
rect 4543 2302 4558 2336
rect 4698 2302 4713 2336
rect 4747 2302 4849 2336
rect 4407 2268 4558 2302
rect 4698 2268 4849 2302
rect 4407 2234 4509 2268
rect 4543 2234 4558 2268
rect 4698 2234 4713 2268
rect 4747 2234 4849 2268
rect 4407 2200 4558 2234
rect 4698 2200 4849 2234
rect 4407 2166 4509 2200
rect 4543 2166 4558 2200
rect 4698 2166 4713 2200
rect 4747 2166 4849 2200
rect 4407 2132 4558 2166
rect 4698 2132 4849 2166
rect 4407 2098 4509 2132
rect 4543 2098 4558 2132
rect 4698 2098 4713 2132
rect 4747 2098 4849 2132
rect 4407 2064 4558 2098
rect 4698 2064 4849 2098
rect 4407 2030 4509 2064
rect 4543 2030 4558 2064
rect 4698 2030 4713 2064
rect 4747 2030 4849 2064
rect 4407 1996 4558 2030
rect 4698 1996 4849 2030
rect 4407 1962 4509 1996
rect 4543 1962 4558 1996
rect 4698 1962 4713 1996
rect 4747 1962 4849 1996
rect 4407 1928 4558 1962
rect 4698 1928 4849 1962
rect 4407 1894 4509 1928
rect 4543 1894 4558 1928
rect 4698 1894 4713 1928
rect 4747 1894 4849 1928
rect 4407 1860 4558 1894
rect 4698 1860 4849 1894
rect 4407 1826 4509 1860
rect 4543 1826 4558 1860
rect 4698 1826 4713 1860
rect 4747 1826 4849 1860
rect 4407 1792 4558 1826
rect 4698 1792 4849 1826
rect 4407 1758 4509 1792
rect 4543 1758 4558 1792
rect 4698 1758 4713 1792
rect 4747 1758 4849 1792
rect 4407 1724 4558 1758
rect 4698 1724 4849 1758
rect 4407 1690 4509 1724
rect 4543 1690 4558 1724
rect 4698 1690 4713 1724
rect 4747 1690 4849 1724
rect 4407 1656 4558 1690
rect 4698 1656 4849 1690
rect 4407 1622 4509 1656
rect 4543 1622 4558 1656
rect 4698 1622 4713 1656
rect 4747 1622 4849 1656
rect 4407 1552 4558 1622
rect 4698 1552 4849 1622
rect 4969 2482 5279 2552
rect 4969 2448 5071 2482
rect 5105 2448 5143 2482
rect 5177 2448 5279 2482
rect 4969 2414 5279 2448
rect 4969 2380 5071 2414
rect 5105 2380 5143 2414
rect 5177 2380 5279 2414
rect 4969 2346 5279 2380
rect 4969 2312 5071 2346
rect 5105 2312 5143 2346
rect 5177 2312 5279 2346
rect 4969 2278 5279 2312
rect 4969 2244 5071 2278
rect 5105 2244 5143 2278
rect 5177 2244 5279 2278
rect 4969 2210 5279 2244
rect 4969 2176 5071 2210
rect 5105 2176 5143 2210
rect 5177 2176 5279 2210
rect 4969 2142 5279 2176
rect 4969 2108 5071 2142
rect 5105 2108 5143 2142
rect 5177 2108 5279 2142
rect 4969 2074 5279 2108
rect 4969 2040 5071 2074
rect 5105 2040 5143 2074
rect 5177 2040 5279 2074
rect 4969 2006 5279 2040
rect 4969 1972 5071 2006
rect 5105 1972 5143 2006
rect 5177 1972 5279 2006
rect 4969 1938 5279 1972
rect 4969 1904 5071 1938
rect 5105 1904 5143 1938
rect 5177 1904 5279 1938
rect 4969 1870 5279 1904
rect 4969 1836 5071 1870
rect 5105 1836 5143 1870
rect 5177 1836 5279 1870
rect 4969 1802 5279 1836
rect 4969 1768 5071 1802
rect 5105 1768 5143 1802
rect 5177 1768 5279 1802
rect 4969 1734 5279 1768
rect 4969 1700 5071 1734
rect 5105 1700 5143 1734
rect 5177 1700 5279 1734
rect 4969 1666 5279 1700
rect 4969 1632 5071 1666
rect 5105 1632 5143 1666
rect 5177 1632 5279 1666
rect 4969 1598 5279 1632
rect 4969 1564 5071 1598
rect 5105 1564 5143 1598
rect 5177 1564 5279 1598
rect 4969 1552 5279 1564
rect 5399 2540 5550 2552
rect 5690 2540 5841 2552
rect 5399 2506 5501 2540
rect 5535 2506 5550 2540
rect 5690 2506 5705 2540
rect 5739 2506 5841 2540
rect 5399 2472 5550 2506
rect 5690 2472 5841 2506
rect 5399 2438 5501 2472
rect 5535 2438 5550 2472
rect 5690 2438 5705 2472
rect 5739 2438 5841 2472
rect 5399 2404 5550 2438
rect 5690 2404 5841 2438
rect 5399 2370 5501 2404
rect 5535 2370 5550 2404
rect 5690 2370 5705 2404
rect 5739 2370 5841 2404
rect 5399 2336 5550 2370
rect 5690 2336 5841 2370
rect 5399 2302 5501 2336
rect 5535 2302 5550 2336
rect 5690 2302 5705 2336
rect 5739 2302 5841 2336
rect 5399 2268 5550 2302
rect 5690 2268 5841 2302
rect 5399 2234 5501 2268
rect 5535 2234 5550 2268
rect 5690 2234 5705 2268
rect 5739 2234 5841 2268
rect 5399 2200 5550 2234
rect 5690 2200 5841 2234
rect 5399 2166 5501 2200
rect 5535 2166 5550 2200
rect 5690 2166 5705 2200
rect 5739 2166 5841 2200
rect 5399 2132 5550 2166
rect 5690 2132 5841 2166
rect 5399 2098 5501 2132
rect 5535 2098 5550 2132
rect 5690 2098 5705 2132
rect 5739 2098 5841 2132
rect 5399 2064 5550 2098
rect 5690 2064 5841 2098
rect 5399 2030 5501 2064
rect 5535 2030 5550 2064
rect 5690 2030 5705 2064
rect 5739 2030 5841 2064
rect 5399 1996 5550 2030
rect 5690 1996 5841 2030
rect 5399 1962 5501 1996
rect 5535 1962 5550 1996
rect 5690 1962 5705 1996
rect 5739 1962 5841 1996
rect 5399 1928 5550 1962
rect 5690 1928 5841 1962
rect 5399 1894 5501 1928
rect 5535 1894 5550 1928
rect 5690 1894 5705 1928
rect 5739 1894 5841 1928
rect 5399 1860 5550 1894
rect 5690 1860 5841 1894
rect 5399 1826 5501 1860
rect 5535 1826 5550 1860
rect 5690 1826 5705 1860
rect 5739 1826 5841 1860
rect 5399 1792 5550 1826
rect 5690 1792 5841 1826
rect 5399 1758 5501 1792
rect 5535 1758 5550 1792
rect 5690 1758 5705 1792
rect 5739 1758 5841 1792
rect 5399 1724 5550 1758
rect 5690 1724 5841 1758
rect 5399 1690 5501 1724
rect 5535 1690 5550 1724
rect 5690 1690 5705 1724
rect 5739 1690 5841 1724
rect 5399 1656 5550 1690
rect 5690 1656 5841 1690
rect 5399 1622 5501 1656
rect 5535 1622 5550 1656
rect 5690 1622 5705 1656
rect 5739 1622 5841 1656
rect 5399 1552 5550 1622
rect 5690 1552 5841 1622
rect 5961 2482 6271 2552
rect 5961 2448 6063 2482
rect 6097 2448 6135 2482
rect 6169 2448 6271 2482
rect 5961 2414 6271 2448
rect 5961 2380 6063 2414
rect 6097 2380 6135 2414
rect 6169 2380 6271 2414
rect 5961 2346 6271 2380
rect 5961 2312 6063 2346
rect 6097 2312 6135 2346
rect 6169 2312 6271 2346
rect 5961 2278 6271 2312
rect 5961 2244 6063 2278
rect 6097 2244 6135 2278
rect 6169 2244 6271 2278
rect 5961 2210 6271 2244
rect 5961 2176 6063 2210
rect 6097 2176 6135 2210
rect 6169 2176 6271 2210
rect 5961 2142 6271 2176
rect 5961 2108 6063 2142
rect 6097 2108 6135 2142
rect 6169 2108 6271 2142
rect 5961 2074 6271 2108
rect 5961 2040 6063 2074
rect 6097 2040 6135 2074
rect 6169 2040 6271 2074
rect 5961 2006 6271 2040
rect 5961 1972 6063 2006
rect 6097 1972 6135 2006
rect 6169 1972 6271 2006
rect 5961 1938 6271 1972
rect 5961 1904 6063 1938
rect 6097 1904 6135 1938
rect 6169 1904 6271 1938
rect 5961 1870 6271 1904
rect 5961 1836 6063 1870
rect 6097 1836 6135 1870
rect 6169 1836 6271 1870
rect 5961 1802 6271 1836
rect 5961 1768 6063 1802
rect 6097 1768 6135 1802
rect 6169 1768 6271 1802
rect 5961 1734 6271 1768
rect 5961 1700 6063 1734
rect 6097 1700 6135 1734
rect 6169 1700 6271 1734
rect 5961 1666 6271 1700
rect 5961 1632 6063 1666
rect 6097 1632 6135 1666
rect 6169 1632 6271 1666
rect 5961 1598 6271 1632
rect 5961 1564 6063 1598
rect 6097 1564 6135 1598
rect 6169 1564 6271 1598
rect 5961 1552 6271 1564
rect 6391 2540 6542 2552
rect 6682 2540 6833 2552
rect 6391 2506 6493 2540
rect 6527 2506 6542 2540
rect 6682 2506 6697 2540
rect 6731 2506 6833 2540
rect 6391 2472 6542 2506
rect 6682 2472 6833 2506
rect 6391 2438 6493 2472
rect 6527 2438 6542 2472
rect 6682 2438 6697 2472
rect 6731 2438 6833 2472
rect 6391 2404 6542 2438
rect 6682 2404 6833 2438
rect 6391 2370 6493 2404
rect 6527 2370 6542 2404
rect 6682 2370 6697 2404
rect 6731 2370 6833 2404
rect 6391 2336 6542 2370
rect 6682 2336 6833 2370
rect 6391 2302 6493 2336
rect 6527 2302 6542 2336
rect 6682 2302 6697 2336
rect 6731 2302 6833 2336
rect 6391 2268 6542 2302
rect 6682 2268 6833 2302
rect 6391 2234 6493 2268
rect 6527 2234 6542 2268
rect 6682 2234 6697 2268
rect 6731 2234 6833 2268
rect 6391 2200 6542 2234
rect 6682 2200 6833 2234
rect 6391 2166 6493 2200
rect 6527 2166 6542 2200
rect 6682 2166 6697 2200
rect 6731 2166 6833 2200
rect 6391 2132 6542 2166
rect 6682 2132 6833 2166
rect 6391 2098 6493 2132
rect 6527 2098 6542 2132
rect 6682 2098 6697 2132
rect 6731 2098 6833 2132
rect 6391 2064 6542 2098
rect 6682 2064 6833 2098
rect 6391 2030 6493 2064
rect 6527 2030 6542 2064
rect 6682 2030 6697 2064
rect 6731 2030 6833 2064
rect 6391 1996 6542 2030
rect 6682 1996 6833 2030
rect 6391 1962 6493 1996
rect 6527 1962 6542 1996
rect 6682 1962 6697 1996
rect 6731 1962 6833 1996
rect 6391 1928 6542 1962
rect 6682 1928 6833 1962
rect 6391 1894 6493 1928
rect 6527 1894 6542 1928
rect 6682 1894 6697 1928
rect 6731 1894 6833 1928
rect 6391 1860 6542 1894
rect 6682 1860 6833 1894
rect 6391 1826 6493 1860
rect 6527 1826 6542 1860
rect 6682 1826 6697 1860
rect 6731 1826 6833 1860
rect 6391 1792 6542 1826
rect 6682 1792 6833 1826
rect 6391 1758 6493 1792
rect 6527 1758 6542 1792
rect 6682 1758 6697 1792
rect 6731 1758 6833 1792
rect 6391 1724 6542 1758
rect 6682 1724 6833 1758
rect 6391 1690 6493 1724
rect 6527 1690 6542 1724
rect 6682 1690 6697 1724
rect 6731 1690 6833 1724
rect 6391 1656 6542 1690
rect 6682 1656 6833 1690
rect 6391 1622 6493 1656
rect 6527 1622 6542 1656
rect 6682 1622 6697 1656
rect 6731 1622 6833 1656
rect 6391 1552 6542 1622
rect 6682 1552 6833 1622
rect 6953 2482 7263 2552
rect 6953 2448 7055 2482
rect 7089 2448 7127 2482
rect 7161 2448 7263 2482
rect 6953 2414 7263 2448
rect 6953 2380 7055 2414
rect 7089 2380 7127 2414
rect 7161 2380 7263 2414
rect 6953 2346 7263 2380
rect 6953 2312 7055 2346
rect 7089 2312 7127 2346
rect 7161 2312 7263 2346
rect 6953 2278 7263 2312
rect 6953 2244 7055 2278
rect 7089 2244 7127 2278
rect 7161 2244 7263 2278
rect 6953 2210 7263 2244
rect 6953 2176 7055 2210
rect 7089 2176 7127 2210
rect 7161 2176 7263 2210
rect 6953 2142 7263 2176
rect 6953 2108 7055 2142
rect 7089 2108 7127 2142
rect 7161 2108 7263 2142
rect 6953 2074 7263 2108
rect 6953 2040 7055 2074
rect 7089 2040 7127 2074
rect 7161 2040 7263 2074
rect 6953 2006 7263 2040
rect 6953 1972 7055 2006
rect 7089 1972 7127 2006
rect 7161 1972 7263 2006
rect 6953 1938 7263 1972
rect 6953 1904 7055 1938
rect 7089 1904 7127 1938
rect 7161 1904 7263 1938
rect 6953 1870 7263 1904
rect 6953 1836 7055 1870
rect 7089 1836 7127 1870
rect 7161 1836 7263 1870
rect 6953 1802 7263 1836
rect 6953 1768 7055 1802
rect 7089 1768 7127 1802
rect 7161 1768 7263 1802
rect 6953 1734 7263 1768
rect 6953 1700 7055 1734
rect 7089 1700 7127 1734
rect 7161 1700 7263 1734
rect 6953 1666 7263 1700
rect 6953 1632 7055 1666
rect 7089 1632 7127 1666
rect 7161 1632 7263 1666
rect 6953 1598 7263 1632
rect 6953 1564 7055 1598
rect 7089 1564 7127 1598
rect 7161 1564 7263 1598
rect 6953 1552 7263 1564
rect 7383 2540 7534 2552
rect 7674 2540 7825 2552
rect 7383 2506 7485 2540
rect 7519 2506 7534 2540
rect 7674 2506 7689 2540
rect 7723 2506 7825 2540
rect 7383 2472 7534 2506
rect 7674 2472 7825 2506
rect 7383 2438 7485 2472
rect 7519 2438 7534 2472
rect 7674 2438 7689 2472
rect 7723 2438 7825 2472
rect 7383 2404 7534 2438
rect 7674 2404 7825 2438
rect 7383 2370 7485 2404
rect 7519 2370 7534 2404
rect 7674 2370 7689 2404
rect 7723 2370 7825 2404
rect 7383 2336 7534 2370
rect 7674 2336 7825 2370
rect 7383 2302 7485 2336
rect 7519 2302 7534 2336
rect 7674 2302 7689 2336
rect 7723 2302 7825 2336
rect 7383 2268 7534 2302
rect 7674 2268 7825 2302
rect 7383 2234 7485 2268
rect 7519 2234 7534 2268
rect 7674 2234 7689 2268
rect 7723 2234 7825 2268
rect 7383 2200 7534 2234
rect 7674 2200 7825 2234
rect 7383 2166 7485 2200
rect 7519 2166 7534 2200
rect 7674 2166 7689 2200
rect 7723 2166 7825 2200
rect 7383 2132 7534 2166
rect 7674 2132 7825 2166
rect 7383 2098 7485 2132
rect 7519 2098 7534 2132
rect 7674 2098 7689 2132
rect 7723 2098 7825 2132
rect 7383 2064 7534 2098
rect 7674 2064 7825 2098
rect 7383 2030 7485 2064
rect 7519 2030 7534 2064
rect 7674 2030 7689 2064
rect 7723 2030 7825 2064
rect 7383 1996 7534 2030
rect 7674 1996 7825 2030
rect 7383 1962 7485 1996
rect 7519 1962 7534 1996
rect 7674 1962 7689 1996
rect 7723 1962 7825 1996
rect 7383 1928 7534 1962
rect 7674 1928 7825 1962
rect 7383 1894 7485 1928
rect 7519 1894 7534 1928
rect 7674 1894 7689 1928
rect 7723 1894 7825 1928
rect 7383 1860 7534 1894
rect 7674 1860 7825 1894
rect 7383 1826 7485 1860
rect 7519 1826 7534 1860
rect 7674 1826 7689 1860
rect 7723 1826 7825 1860
rect 7383 1792 7534 1826
rect 7674 1792 7825 1826
rect 7383 1758 7485 1792
rect 7519 1758 7534 1792
rect 7674 1758 7689 1792
rect 7723 1758 7825 1792
rect 7383 1724 7534 1758
rect 7674 1724 7825 1758
rect 7383 1690 7485 1724
rect 7519 1690 7534 1724
rect 7674 1690 7689 1724
rect 7723 1690 7825 1724
rect 7383 1656 7534 1690
rect 7674 1656 7825 1690
rect 7383 1622 7485 1656
rect 7519 1622 7534 1656
rect 7674 1622 7689 1656
rect 7723 1622 7825 1656
rect 7383 1552 7534 1622
rect 7674 1552 7825 1622
rect 7945 2482 8255 2552
rect 7945 2448 8047 2482
rect 8081 2448 8119 2482
rect 8153 2448 8255 2482
rect 7945 2414 8255 2448
rect 7945 2380 8047 2414
rect 8081 2380 8119 2414
rect 8153 2380 8255 2414
rect 7945 2346 8255 2380
rect 7945 2312 8047 2346
rect 8081 2312 8119 2346
rect 8153 2312 8255 2346
rect 7945 2278 8255 2312
rect 7945 2244 8047 2278
rect 8081 2244 8119 2278
rect 8153 2244 8255 2278
rect 7945 2210 8255 2244
rect 7945 2176 8047 2210
rect 8081 2176 8119 2210
rect 8153 2176 8255 2210
rect 7945 2142 8255 2176
rect 7945 2108 8047 2142
rect 8081 2108 8119 2142
rect 8153 2108 8255 2142
rect 7945 2074 8255 2108
rect 7945 2040 8047 2074
rect 8081 2040 8119 2074
rect 8153 2040 8255 2074
rect 7945 2006 8255 2040
rect 7945 1972 8047 2006
rect 8081 1972 8119 2006
rect 8153 1972 8255 2006
rect 7945 1938 8255 1972
rect 7945 1904 8047 1938
rect 8081 1904 8119 1938
rect 8153 1904 8255 1938
rect 7945 1870 8255 1904
rect 7945 1836 8047 1870
rect 8081 1836 8119 1870
rect 8153 1836 8255 1870
rect 7945 1802 8255 1836
rect 7945 1768 8047 1802
rect 8081 1768 8119 1802
rect 8153 1768 8255 1802
rect 7945 1734 8255 1768
rect 7945 1700 8047 1734
rect 8081 1700 8119 1734
rect 8153 1700 8255 1734
rect 7945 1666 8255 1700
rect 7945 1632 8047 1666
rect 8081 1632 8119 1666
rect 8153 1632 8255 1666
rect 7945 1598 8255 1632
rect 7945 1564 8047 1598
rect 8081 1564 8119 1598
rect 8153 1564 8255 1598
rect 7945 1552 8255 1564
rect 8375 2540 8526 2552
rect 8666 2540 8817 2552
rect 8375 2506 8477 2540
rect 8511 2506 8526 2540
rect 8666 2506 8681 2540
rect 8715 2506 8817 2540
rect 8375 2472 8526 2506
rect 8666 2472 8817 2506
rect 8375 2438 8477 2472
rect 8511 2438 8526 2472
rect 8666 2438 8681 2472
rect 8715 2438 8817 2472
rect 8375 2404 8526 2438
rect 8666 2404 8817 2438
rect 8375 2370 8477 2404
rect 8511 2370 8526 2404
rect 8666 2370 8681 2404
rect 8715 2370 8817 2404
rect 8375 2336 8526 2370
rect 8666 2336 8817 2370
rect 8375 2302 8477 2336
rect 8511 2302 8526 2336
rect 8666 2302 8681 2336
rect 8715 2302 8817 2336
rect 8375 2268 8526 2302
rect 8666 2268 8817 2302
rect 8375 2234 8477 2268
rect 8511 2234 8526 2268
rect 8666 2234 8681 2268
rect 8715 2234 8817 2268
rect 8375 2200 8526 2234
rect 8666 2200 8817 2234
rect 8375 2166 8477 2200
rect 8511 2166 8526 2200
rect 8666 2166 8681 2200
rect 8715 2166 8817 2200
rect 8375 2132 8526 2166
rect 8666 2132 8817 2166
rect 8375 2098 8477 2132
rect 8511 2098 8526 2132
rect 8666 2098 8681 2132
rect 8715 2098 8817 2132
rect 8375 2064 8526 2098
rect 8666 2064 8817 2098
rect 8375 2030 8477 2064
rect 8511 2030 8526 2064
rect 8666 2030 8681 2064
rect 8715 2030 8817 2064
rect 8375 1996 8526 2030
rect 8666 1996 8817 2030
rect 8375 1962 8477 1996
rect 8511 1962 8526 1996
rect 8666 1962 8681 1996
rect 8715 1962 8817 1996
rect 8375 1928 8526 1962
rect 8666 1928 8817 1962
rect 8375 1894 8477 1928
rect 8511 1894 8526 1928
rect 8666 1894 8681 1928
rect 8715 1894 8817 1928
rect 8375 1860 8526 1894
rect 8666 1860 8817 1894
rect 8375 1826 8477 1860
rect 8511 1826 8526 1860
rect 8666 1826 8681 1860
rect 8715 1826 8817 1860
rect 8375 1792 8526 1826
rect 8666 1792 8817 1826
rect 8375 1758 8477 1792
rect 8511 1758 8526 1792
rect 8666 1758 8681 1792
rect 8715 1758 8817 1792
rect 8375 1724 8526 1758
rect 8666 1724 8817 1758
rect 8375 1690 8477 1724
rect 8511 1690 8526 1724
rect 8666 1690 8681 1724
rect 8715 1690 8817 1724
rect 8375 1656 8526 1690
rect 8666 1656 8817 1690
rect 8375 1622 8477 1656
rect 8511 1622 8526 1656
rect 8666 1622 8681 1656
rect 8715 1622 8817 1656
rect 8375 1552 8526 1622
rect 8666 1552 8817 1622
rect 8937 2482 9247 2552
rect 8937 2448 9039 2482
rect 9073 2448 9111 2482
rect 9145 2448 9247 2482
rect 8937 2414 9247 2448
rect 8937 2380 9039 2414
rect 9073 2380 9111 2414
rect 9145 2380 9247 2414
rect 8937 2346 9247 2380
rect 8937 2312 9039 2346
rect 9073 2312 9111 2346
rect 9145 2312 9247 2346
rect 8937 2278 9247 2312
rect 8937 2244 9039 2278
rect 9073 2244 9111 2278
rect 9145 2244 9247 2278
rect 8937 2210 9247 2244
rect 8937 2176 9039 2210
rect 9073 2176 9111 2210
rect 9145 2176 9247 2210
rect 8937 2142 9247 2176
rect 8937 2108 9039 2142
rect 9073 2108 9111 2142
rect 9145 2108 9247 2142
rect 8937 2074 9247 2108
rect 8937 2040 9039 2074
rect 9073 2040 9111 2074
rect 9145 2040 9247 2074
rect 8937 2006 9247 2040
rect 8937 1972 9039 2006
rect 9073 1972 9111 2006
rect 9145 1972 9247 2006
rect 8937 1938 9247 1972
rect 8937 1904 9039 1938
rect 9073 1904 9111 1938
rect 9145 1904 9247 1938
rect 8937 1870 9247 1904
rect 8937 1836 9039 1870
rect 9073 1836 9111 1870
rect 9145 1836 9247 1870
rect 8937 1802 9247 1836
rect 8937 1768 9039 1802
rect 9073 1768 9111 1802
rect 9145 1768 9247 1802
rect 8937 1734 9247 1768
rect 8937 1700 9039 1734
rect 9073 1700 9111 1734
rect 9145 1700 9247 1734
rect 8937 1666 9247 1700
rect 8937 1632 9039 1666
rect 9073 1632 9111 1666
rect 9145 1632 9247 1666
rect 8937 1598 9247 1632
rect 8937 1564 9039 1598
rect 9073 1564 9111 1598
rect 9145 1564 9247 1598
rect 8937 1552 9247 1564
rect 9367 2540 9518 2552
rect 9658 2540 9809 2552
rect 9367 2506 9469 2540
rect 9503 2506 9518 2540
rect 9658 2506 9673 2540
rect 9707 2506 9809 2540
rect 9367 2472 9518 2506
rect 9658 2472 9809 2506
rect 9367 2438 9469 2472
rect 9503 2438 9518 2472
rect 9658 2438 9673 2472
rect 9707 2438 9809 2472
rect 9367 2404 9518 2438
rect 9658 2404 9809 2438
rect 9367 2370 9469 2404
rect 9503 2370 9518 2404
rect 9658 2370 9673 2404
rect 9707 2370 9809 2404
rect 9367 2336 9518 2370
rect 9658 2336 9809 2370
rect 9367 2302 9469 2336
rect 9503 2302 9518 2336
rect 9658 2302 9673 2336
rect 9707 2302 9809 2336
rect 9367 2268 9518 2302
rect 9658 2268 9809 2302
rect 9367 2234 9469 2268
rect 9503 2234 9518 2268
rect 9658 2234 9673 2268
rect 9707 2234 9809 2268
rect 9367 2200 9518 2234
rect 9658 2200 9809 2234
rect 9367 2166 9469 2200
rect 9503 2166 9518 2200
rect 9658 2166 9673 2200
rect 9707 2166 9809 2200
rect 9367 2132 9518 2166
rect 9658 2132 9809 2166
rect 9367 2098 9469 2132
rect 9503 2098 9518 2132
rect 9658 2098 9673 2132
rect 9707 2098 9809 2132
rect 9367 2064 9518 2098
rect 9658 2064 9809 2098
rect 9367 2030 9469 2064
rect 9503 2030 9518 2064
rect 9658 2030 9673 2064
rect 9707 2030 9809 2064
rect 9367 1996 9518 2030
rect 9658 1996 9809 2030
rect 9367 1962 9469 1996
rect 9503 1962 9518 1996
rect 9658 1962 9673 1996
rect 9707 1962 9809 1996
rect 9367 1928 9518 1962
rect 9658 1928 9809 1962
rect 9367 1894 9469 1928
rect 9503 1894 9518 1928
rect 9658 1894 9673 1928
rect 9707 1894 9809 1928
rect 9367 1860 9518 1894
rect 9658 1860 9809 1894
rect 9367 1826 9469 1860
rect 9503 1826 9518 1860
rect 9658 1826 9673 1860
rect 9707 1826 9809 1860
rect 9367 1792 9518 1826
rect 9658 1792 9809 1826
rect 9367 1758 9469 1792
rect 9503 1758 9518 1792
rect 9658 1758 9673 1792
rect 9707 1758 9809 1792
rect 9367 1724 9518 1758
rect 9658 1724 9809 1758
rect 9367 1690 9469 1724
rect 9503 1690 9518 1724
rect 9658 1690 9673 1724
rect 9707 1690 9809 1724
rect 9367 1656 9518 1690
rect 9658 1656 9809 1690
rect 9367 1622 9469 1656
rect 9503 1622 9518 1656
rect 9658 1622 9673 1656
rect 9707 1622 9809 1656
rect 9367 1552 9518 1622
rect 9658 1552 9809 1622
rect 9929 2482 10239 2552
rect 9929 2448 10031 2482
rect 10065 2448 10103 2482
rect 10137 2448 10239 2482
rect 9929 2414 10239 2448
rect 9929 2380 10031 2414
rect 10065 2380 10103 2414
rect 10137 2380 10239 2414
rect 9929 2346 10239 2380
rect 9929 2312 10031 2346
rect 10065 2312 10103 2346
rect 10137 2312 10239 2346
rect 9929 2278 10239 2312
rect 9929 2244 10031 2278
rect 10065 2244 10103 2278
rect 10137 2244 10239 2278
rect 9929 2210 10239 2244
rect 9929 2176 10031 2210
rect 10065 2176 10103 2210
rect 10137 2176 10239 2210
rect 9929 2142 10239 2176
rect 9929 2108 10031 2142
rect 10065 2108 10103 2142
rect 10137 2108 10239 2142
rect 9929 2074 10239 2108
rect 9929 2040 10031 2074
rect 10065 2040 10103 2074
rect 10137 2040 10239 2074
rect 9929 2006 10239 2040
rect 9929 1972 10031 2006
rect 10065 1972 10103 2006
rect 10137 1972 10239 2006
rect 9929 1938 10239 1972
rect 9929 1904 10031 1938
rect 10065 1904 10103 1938
rect 10137 1904 10239 1938
rect 9929 1870 10239 1904
rect 9929 1836 10031 1870
rect 10065 1836 10103 1870
rect 10137 1836 10239 1870
rect 9929 1802 10239 1836
rect 9929 1768 10031 1802
rect 10065 1768 10103 1802
rect 10137 1768 10239 1802
rect 9929 1734 10239 1768
rect 9929 1700 10031 1734
rect 10065 1700 10103 1734
rect 10137 1700 10239 1734
rect 9929 1666 10239 1700
rect 9929 1632 10031 1666
rect 10065 1632 10103 1666
rect 10137 1632 10239 1666
rect 9929 1598 10239 1632
rect 9929 1564 10031 1598
rect 10065 1564 10103 1598
rect 10137 1564 10239 1598
rect 9929 1552 10239 1564
rect 10359 2540 10510 2552
rect 10650 2540 10801 2552
rect 10359 2506 10461 2540
rect 10495 2506 10510 2540
rect 10650 2506 10665 2540
rect 10699 2506 10801 2540
rect 10359 2472 10510 2506
rect 10650 2472 10801 2506
rect 10359 2438 10461 2472
rect 10495 2438 10510 2472
rect 10650 2438 10665 2472
rect 10699 2438 10801 2472
rect 10359 2404 10510 2438
rect 10650 2404 10801 2438
rect 10359 2370 10461 2404
rect 10495 2370 10510 2404
rect 10650 2370 10665 2404
rect 10699 2370 10801 2404
rect 10359 2336 10510 2370
rect 10650 2336 10801 2370
rect 10359 2302 10461 2336
rect 10495 2302 10510 2336
rect 10650 2302 10665 2336
rect 10699 2302 10801 2336
rect 10359 2268 10510 2302
rect 10650 2268 10801 2302
rect 10359 2234 10461 2268
rect 10495 2234 10510 2268
rect 10650 2234 10665 2268
rect 10699 2234 10801 2268
rect 10359 2200 10510 2234
rect 10650 2200 10801 2234
rect 10359 2166 10461 2200
rect 10495 2166 10510 2200
rect 10650 2166 10665 2200
rect 10699 2166 10801 2200
rect 10359 2132 10510 2166
rect 10650 2132 10801 2166
rect 10359 2098 10461 2132
rect 10495 2098 10510 2132
rect 10650 2098 10665 2132
rect 10699 2098 10801 2132
rect 10359 2064 10510 2098
rect 10650 2064 10801 2098
rect 10359 2030 10461 2064
rect 10495 2030 10510 2064
rect 10650 2030 10665 2064
rect 10699 2030 10801 2064
rect 10359 1996 10510 2030
rect 10650 1996 10801 2030
rect 10359 1962 10461 1996
rect 10495 1962 10510 1996
rect 10650 1962 10665 1996
rect 10699 1962 10801 1996
rect 10359 1928 10510 1962
rect 10650 1928 10801 1962
rect 10359 1894 10461 1928
rect 10495 1894 10510 1928
rect 10650 1894 10665 1928
rect 10699 1894 10801 1928
rect 10359 1860 10510 1894
rect 10650 1860 10801 1894
rect 10359 1826 10461 1860
rect 10495 1826 10510 1860
rect 10650 1826 10665 1860
rect 10699 1826 10801 1860
rect 10359 1792 10510 1826
rect 10650 1792 10801 1826
rect 10359 1758 10461 1792
rect 10495 1758 10510 1792
rect 10650 1758 10665 1792
rect 10699 1758 10801 1792
rect 10359 1724 10510 1758
rect 10650 1724 10801 1758
rect 10359 1690 10461 1724
rect 10495 1690 10510 1724
rect 10650 1690 10665 1724
rect 10699 1690 10801 1724
rect 10359 1656 10510 1690
rect 10650 1656 10801 1690
rect 10359 1622 10461 1656
rect 10495 1622 10510 1656
rect 10650 1622 10665 1656
rect 10699 1622 10801 1656
rect 10359 1552 10510 1622
rect 10650 1552 10801 1622
rect 10921 2482 11231 2552
rect 10921 2448 11023 2482
rect 11057 2448 11095 2482
rect 11129 2448 11231 2482
rect 10921 2414 11231 2448
rect 10921 2380 11023 2414
rect 11057 2380 11095 2414
rect 11129 2380 11231 2414
rect 10921 2346 11231 2380
rect 10921 2312 11023 2346
rect 11057 2312 11095 2346
rect 11129 2312 11231 2346
rect 10921 2278 11231 2312
rect 10921 2244 11023 2278
rect 11057 2244 11095 2278
rect 11129 2244 11231 2278
rect 10921 2210 11231 2244
rect 10921 2176 11023 2210
rect 11057 2176 11095 2210
rect 11129 2176 11231 2210
rect 10921 2142 11231 2176
rect 10921 2108 11023 2142
rect 11057 2108 11095 2142
rect 11129 2108 11231 2142
rect 10921 2074 11231 2108
rect 10921 2040 11023 2074
rect 11057 2040 11095 2074
rect 11129 2040 11231 2074
rect 10921 2006 11231 2040
rect 10921 1972 11023 2006
rect 11057 1972 11095 2006
rect 11129 1972 11231 2006
rect 10921 1938 11231 1972
rect 10921 1904 11023 1938
rect 11057 1904 11095 1938
rect 11129 1904 11231 1938
rect 10921 1870 11231 1904
rect 10921 1836 11023 1870
rect 11057 1836 11095 1870
rect 11129 1836 11231 1870
rect 10921 1802 11231 1836
rect 10921 1768 11023 1802
rect 11057 1768 11095 1802
rect 11129 1768 11231 1802
rect 10921 1734 11231 1768
rect 10921 1700 11023 1734
rect 11057 1700 11095 1734
rect 11129 1700 11231 1734
rect 10921 1666 11231 1700
rect 10921 1632 11023 1666
rect 11057 1632 11095 1666
rect 11129 1632 11231 1666
rect 10921 1598 11231 1632
rect 10921 1564 11023 1598
rect 11057 1564 11095 1598
rect 11129 1564 11231 1598
rect 10921 1552 11231 1564
rect 11351 2540 11502 2552
rect 11642 2540 11793 2552
rect 11351 2506 11453 2540
rect 11487 2506 11502 2540
rect 11642 2506 11657 2540
rect 11691 2506 11793 2540
rect 11351 2472 11502 2506
rect 11642 2472 11793 2506
rect 11351 2438 11453 2472
rect 11487 2438 11502 2472
rect 11642 2438 11657 2472
rect 11691 2438 11793 2472
rect 11351 2404 11502 2438
rect 11642 2404 11793 2438
rect 11351 2370 11453 2404
rect 11487 2370 11502 2404
rect 11642 2370 11657 2404
rect 11691 2370 11793 2404
rect 11351 2336 11502 2370
rect 11642 2336 11793 2370
rect 11351 2302 11453 2336
rect 11487 2302 11502 2336
rect 11642 2302 11657 2336
rect 11691 2302 11793 2336
rect 11351 2268 11502 2302
rect 11642 2268 11793 2302
rect 11351 2234 11453 2268
rect 11487 2234 11502 2268
rect 11642 2234 11657 2268
rect 11691 2234 11793 2268
rect 11351 2200 11502 2234
rect 11642 2200 11793 2234
rect 11351 2166 11453 2200
rect 11487 2166 11502 2200
rect 11642 2166 11657 2200
rect 11691 2166 11793 2200
rect 11351 2132 11502 2166
rect 11642 2132 11793 2166
rect 11351 2098 11453 2132
rect 11487 2098 11502 2132
rect 11642 2098 11657 2132
rect 11691 2098 11793 2132
rect 11351 2064 11502 2098
rect 11642 2064 11793 2098
rect 11351 2030 11453 2064
rect 11487 2030 11502 2064
rect 11642 2030 11657 2064
rect 11691 2030 11793 2064
rect 11351 1996 11502 2030
rect 11642 1996 11793 2030
rect 11351 1962 11453 1996
rect 11487 1962 11502 1996
rect 11642 1962 11657 1996
rect 11691 1962 11793 1996
rect 11351 1928 11502 1962
rect 11642 1928 11793 1962
rect 11351 1894 11453 1928
rect 11487 1894 11502 1928
rect 11642 1894 11657 1928
rect 11691 1894 11793 1928
rect 11351 1860 11502 1894
rect 11642 1860 11793 1894
rect 11351 1826 11453 1860
rect 11487 1826 11502 1860
rect 11642 1826 11657 1860
rect 11691 1826 11793 1860
rect 11351 1792 11502 1826
rect 11642 1792 11793 1826
rect 11351 1758 11453 1792
rect 11487 1758 11502 1792
rect 11642 1758 11657 1792
rect 11691 1758 11793 1792
rect 11351 1724 11502 1758
rect 11642 1724 11793 1758
rect 11351 1690 11453 1724
rect 11487 1690 11502 1724
rect 11642 1690 11657 1724
rect 11691 1690 11793 1724
rect 11351 1656 11502 1690
rect 11642 1656 11793 1690
rect 11351 1622 11453 1656
rect 11487 1622 11502 1656
rect 11642 1622 11657 1656
rect 11691 1622 11793 1656
rect 11351 1552 11502 1622
rect 11642 1552 11793 1622
rect 11913 2482 12223 2552
rect 11913 2448 12015 2482
rect 12049 2448 12087 2482
rect 12121 2448 12223 2482
rect 11913 2414 12223 2448
rect 11913 2380 12015 2414
rect 12049 2380 12087 2414
rect 12121 2380 12223 2414
rect 11913 2346 12223 2380
rect 11913 2312 12015 2346
rect 12049 2312 12087 2346
rect 12121 2312 12223 2346
rect 11913 2278 12223 2312
rect 11913 2244 12015 2278
rect 12049 2244 12087 2278
rect 12121 2244 12223 2278
rect 11913 2210 12223 2244
rect 11913 2176 12015 2210
rect 12049 2176 12087 2210
rect 12121 2176 12223 2210
rect 11913 2142 12223 2176
rect 11913 2108 12015 2142
rect 12049 2108 12087 2142
rect 12121 2108 12223 2142
rect 11913 2074 12223 2108
rect 11913 2040 12015 2074
rect 12049 2040 12087 2074
rect 12121 2040 12223 2074
rect 11913 2006 12223 2040
rect 11913 1972 12015 2006
rect 12049 1972 12087 2006
rect 12121 1972 12223 2006
rect 11913 1938 12223 1972
rect 11913 1904 12015 1938
rect 12049 1904 12087 1938
rect 12121 1904 12223 1938
rect 11913 1870 12223 1904
rect 11913 1836 12015 1870
rect 12049 1836 12087 1870
rect 12121 1836 12223 1870
rect 11913 1802 12223 1836
rect 11913 1768 12015 1802
rect 12049 1768 12087 1802
rect 12121 1768 12223 1802
rect 11913 1734 12223 1768
rect 11913 1700 12015 1734
rect 12049 1700 12087 1734
rect 12121 1700 12223 1734
rect 11913 1666 12223 1700
rect 11913 1632 12015 1666
rect 12049 1632 12087 1666
rect 12121 1632 12223 1666
rect 11913 1598 12223 1632
rect 11913 1564 12015 1598
rect 12049 1564 12087 1598
rect 12121 1564 12223 1598
rect 11913 1552 12223 1564
rect 12343 2540 12494 2552
rect 12634 2540 12785 2552
rect 12343 2506 12445 2540
rect 12479 2506 12494 2540
rect 12634 2506 12649 2540
rect 12683 2506 12785 2540
rect 12343 2472 12494 2506
rect 12634 2472 12785 2506
rect 12343 2438 12445 2472
rect 12479 2438 12494 2472
rect 12634 2438 12649 2472
rect 12683 2438 12785 2472
rect 12343 2404 12494 2438
rect 12634 2404 12785 2438
rect 12343 2370 12445 2404
rect 12479 2370 12494 2404
rect 12634 2370 12649 2404
rect 12683 2370 12785 2404
rect 12343 2336 12494 2370
rect 12634 2336 12785 2370
rect 12343 2302 12445 2336
rect 12479 2302 12494 2336
rect 12634 2302 12649 2336
rect 12683 2302 12785 2336
rect 12343 2268 12494 2302
rect 12634 2268 12785 2302
rect 12343 2234 12445 2268
rect 12479 2234 12494 2268
rect 12634 2234 12649 2268
rect 12683 2234 12785 2268
rect 12343 2200 12494 2234
rect 12634 2200 12785 2234
rect 12343 2166 12445 2200
rect 12479 2166 12494 2200
rect 12634 2166 12649 2200
rect 12683 2166 12785 2200
rect 12343 2132 12494 2166
rect 12634 2132 12785 2166
rect 12343 2098 12445 2132
rect 12479 2098 12494 2132
rect 12634 2098 12649 2132
rect 12683 2098 12785 2132
rect 12343 2064 12494 2098
rect 12634 2064 12785 2098
rect 12343 2030 12445 2064
rect 12479 2030 12494 2064
rect 12634 2030 12649 2064
rect 12683 2030 12785 2064
rect 12343 1996 12494 2030
rect 12634 1996 12785 2030
rect 12343 1962 12445 1996
rect 12479 1962 12494 1996
rect 12634 1962 12649 1996
rect 12683 1962 12785 1996
rect 12343 1928 12494 1962
rect 12634 1928 12785 1962
rect 12343 1894 12445 1928
rect 12479 1894 12494 1928
rect 12634 1894 12649 1928
rect 12683 1894 12785 1928
rect 12343 1860 12494 1894
rect 12634 1860 12785 1894
rect 12343 1826 12445 1860
rect 12479 1826 12494 1860
rect 12634 1826 12649 1860
rect 12683 1826 12785 1860
rect 12343 1792 12494 1826
rect 12634 1792 12785 1826
rect 12343 1758 12445 1792
rect 12479 1758 12494 1792
rect 12634 1758 12649 1792
rect 12683 1758 12785 1792
rect 12343 1724 12494 1758
rect 12634 1724 12785 1758
rect 12343 1690 12445 1724
rect 12479 1690 12494 1724
rect 12634 1690 12649 1724
rect 12683 1690 12785 1724
rect 12343 1656 12494 1690
rect 12634 1656 12785 1690
rect 12343 1622 12445 1656
rect 12479 1622 12494 1656
rect 12634 1622 12649 1656
rect 12683 1622 12785 1656
rect 12343 1552 12494 1622
rect 12634 1552 12785 1622
rect 12905 2482 13215 2552
rect 12905 2448 13007 2482
rect 13041 2448 13079 2482
rect 13113 2448 13215 2482
rect 12905 2414 13215 2448
rect 12905 2380 13007 2414
rect 13041 2380 13079 2414
rect 13113 2380 13215 2414
rect 12905 2346 13215 2380
rect 12905 2312 13007 2346
rect 13041 2312 13079 2346
rect 13113 2312 13215 2346
rect 12905 2278 13215 2312
rect 12905 2244 13007 2278
rect 13041 2244 13079 2278
rect 13113 2244 13215 2278
rect 12905 2210 13215 2244
rect 12905 2176 13007 2210
rect 13041 2176 13079 2210
rect 13113 2176 13215 2210
rect 12905 2142 13215 2176
rect 12905 2108 13007 2142
rect 13041 2108 13079 2142
rect 13113 2108 13215 2142
rect 12905 2074 13215 2108
rect 12905 2040 13007 2074
rect 13041 2040 13079 2074
rect 13113 2040 13215 2074
rect 12905 2006 13215 2040
rect 12905 1972 13007 2006
rect 13041 1972 13079 2006
rect 13113 1972 13215 2006
rect 12905 1938 13215 1972
rect 12905 1904 13007 1938
rect 13041 1904 13079 1938
rect 13113 1904 13215 1938
rect 12905 1870 13215 1904
rect 12905 1836 13007 1870
rect 13041 1836 13079 1870
rect 13113 1836 13215 1870
rect 12905 1802 13215 1836
rect 12905 1768 13007 1802
rect 13041 1768 13079 1802
rect 13113 1768 13215 1802
rect 12905 1734 13215 1768
rect 12905 1700 13007 1734
rect 13041 1700 13079 1734
rect 13113 1700 13215 1734
rect 12905 1666 13215 1700
rect 12905 1632 13007 1666
rect 13041 1632 13079 1666
rect 13113 1632 13215 1666
rect 12905 1598 13215 1632
rect 12905 1564 13007 1598
rect 13041 1564 13079 1598
rect 13113 1564 13215 1598
rect 12905 1552 13215 1564
rect 13335 2540 13486 2552
rect 13626 2540 13777 2552
rect 13335 2506 13437 2540
rect 13471 2506 13486 2540
rect 13626 2506 13641 2540
rect 13675 2506 13777 2540
rect 13335 2472 13486 2506
rect 13626 2472 13777 2506
rect 13335 2438 13437 2472
rect 13471 2438 13486 2472
rect 13626 2438 13641 2472
rect 13675 2438 13777 2472
rect 13335 2404 13486 2438
rect 13626 2404 13777 2438
rect 13335 2370 13437 2404
rect 13471 2370 13486 2404
rect 13626 2370 13641 2404
rect 13675 2370 13777 2404
rect 13335 2336 13486 2370
rect 13626 2336 13777 2370
rect 13335 2302 13437 2336
rect 13471 2302 13486 2336
rect 13626 2302 13641 2336
rect 13675 2302 13777 2336
rect 13335 2268 13486 2302
rect 13626 2268 13777 2302
rect 13335 2234 13437 2268
rect 13471 2234 13486 2268
rect 13626 2234 13641 2268
rect 13675 2234 13777 2268
rect 13335 2200 13486 2234
rect 13626 2200 13777 2234
rect 13335 2166 13437 2200
rect 13471 2166 13486 2200
rect 13626 2166 13641 2200
rect 13675 2166 13777 2200
rect 13335 2132 13486 2166
rect 13626 2132 13777 2166
rect 13335 2098 13437 2132
rect 13471 2098 13486 2132
rect 13626 2098 13641 2132
rect 13675 2098 13777 2132
rect 13335 2064 13486 2098
rect 13626 2064 13777 2098
rect 13335 2030 13437 2064
rect 13471 2030 13486 2064
rect 13626 2030 13641 2064
rect 13675 2030 13777 2064
rect 13335 1996 13486 2030
rect 13626 1996 13777 2030
rect 13335 1962 13437 1996
rect 13471 1962 13486 1996
rect 13626 1962 13641 1996
rect 13675 1962 13777 1996
rect 13335 1928 13486 1962
rect 13626 1928 13777 1962
rect 13335 1894 13437 1928
rect 13471 1894 13486 1928
rect 13626 1894 13641 1928
rect 13675 1894 13777 1928
rect 13335 1860 13486 1894
rect 13626 1860 13777 1894
rect 13335 1826 13437 1860
rect 13471 1826 13486 1860
rect 13626 1826 13641 1860
rect 13675 1826 13777 1860
rect 13335 1792 13486 1826
rect 13626 1792 13777 1826
rect 13335 1758 13437 1792
rect 13471 1758 13486 1792
rect 13626 1758 13641 1792
rect 13675 1758 13777 1792
rect 13335 1724 13486 1758
rect 13626 1724 13777 1758
rect 13335 1690 13437 1724
rect 13471 1690 13486 1724
rect 13626 1690 13641 1724
rect 13675 1690 13777 1724
rect 13335 1656 13486 1690
rect 13626 1656 13777 1690
rect 13335 1622 13437 1656
rect 13471 1622 13486 1656
rect 13626 1622 13641 1656
rect 13675 1622 13777 1656
rect 13335 1552 13486 1622
rect 13626 1552 13777 1622
rect 13897 2482 14135 2552
rect 13897 2448 13999 2482
rect 14033 2448 14135 2482
rect 13897 2414 14135 2448
rect 13897 2380 13999 2414
rect 14033 2380 14135 2414
rect 13897 2346 14135 2380
rect 13897 2312 13999 2346
rect 14033 2312 14135 2346
rect 13897 2278 14135 2312
rect 13897 2244 13999 2278
rect 14033 2244 14135 2278
rect 13897 2210 14135 2244
rect 13897 2176 13999 2210
rect 14033 2176 14135 2210
rect 13897 2142 14135 2176
rect 13897 2108 13999 2142
rect 14033 2108 14135 2142
rect 13897 2074 14135 2108
rect 13897 2040 13999 2074
rect 14033 2040 14135 2074
rect 13897 2006 14135 2040
rect 13897 1972 13999 2006
rect 14033 1972 14135 2006
rect 13897 1938 14135 1972
rect 13897 1904 13999 1938
rect 14033 1904 14135 1938
rect 13897 1870 14135 1904
rect 13897 1836 13999 1870
rect 14033 1836 14135 1870
rect 13897 1802 14135 1836
rect 13897 1768 13999 1802
rect 14033 1768 14135 1802
rect 13897 1734 14135 1768
rect 13897 1700 13999 1734
rect 14033 1700 14135 1734
rect 13897 1666 14135 1700
rect 13897 1632 13999 1666
rect 14033 1632 14135 1666
rect 13897 1598 14135 1632
rect 13897 1564 13999 1598
rect 14033 1564 14135 1598
rect 13897 1552 14135 1564
rect 14255 2482 14427 2552
rect 14255 2448 14356 2482
rect 14390 2448 14427 2482
rect 14255 2414 14427 2448
rect 14255 2380 14356 2414
rect 14390 2380 14427 2414
rect 14255 2346 14427 2380
rect 14255 2312 14356 2346
rect 14390 2312 14427 2346
rect 14255 2278 14427 2312
rect 14255 2244 14356 2278
rect 14390 2244 14427 2278
rect 14255 2210 14427 2244
rect 14255 2176 14356 2210
rect 14390 2176 14427 2210
rect 14255 2142 14427 2176
rect 14255 2108 14356 2142
rect 14390 2108 14427 2142
rect 14255 2074 14427 2108
rect 14255 2040 14356 2074
rect 14390 2040 14427 2074
rect 14255 2006 14427 2040
rect 14255 1972 14356 2006
rect 14390 1972 14427 2006
rect 14255 1938 14427 1972
rect 14255 1904 14356 1938
rect 14390 1904 14427 1938
rect 14255 1870 14427 1904
rect 14255 1836 14356 1870
rect 14390 1836 14427 1870
rect 14255 1802 14427 1836
rect 14255 1768 14356 1802
rect 14390 1768 14427 1802
rect 14255 1734 14427 1768
rect 14255 1700 14356 1734
rect 14390 1700 14427 1734
rect 14255 1666 14427 1700
rect 14255 1632 14356 1666
rect 14390 1632 14427 1666
rect 14255 1598 14427 1632
rect 14255 1564 14356 1598
rect 14390 1564 14427 1598
rect 14255 1552 14427 1564
<< mvpdiffc >>
rect 745 4048 779 4082
rect 745 3980 779 4014
rect 745 3912 779 3946
rect 745 3844 779 3878
rect 745 3776 779 3810
rect 745 3708 779 3742
rect 745 3640 779 3674
rect 745 3572 779 3606
rect 745 3504 779 3538
rect 745 3436 779 3470
rect 745 3368 779 3402
rect 745 3300 779 3334
rect 745 3232 779 3266
rect 745 3164 779 3198
rect 1103 4048 1137 4082
rect 1175 4048 1209 4082
rect 1103 3980 1137 4014
rect 1175 3980 1209 4014
rect 1103 3912 1137 3946
rect 1175 3912 1209 3946
rect 1103 3844 1137 3878
rect 1175 3844 1209 3878
rect 1103 3776 1137 3810
rect 1175 3776 1209 3810
rect 1103 3708 1137 3742
rect 1175 3708 1209 3742
rect 1103 3640 1137 3674
rect 1175 3640 1209 3674
rect 1103 3572 1137 3606
rect 1175 3572 1209 3606
rect 1103 3504 1137 3538
rect 1175 3504 1209 3538
rect 1103 3436 1137 3470
rect 1175 3436 1209 3470
rect 1103 3368 1137 3402
rect 1175 3368 1209 3402
rect 1103 3300 1137 3334
rect 1175 3300 1209 3334
rect 1103 3232 1137 3266
rect 1175 3232 1209 3266
rect 1103 3164 1137 3198
rect 1175 3164 1209 3198
rect 1533 4048 1567 4082
rect 1737 4048 1771 4082
rect 1533 3980 1567 4014
rect 1737 3980 1771 4014
rect 1533 3912 1567 3946
rect 1737 3912 1771 3946
rect 1533 3844 1567 3878
rect 1737 3844 1771 3878
rect 1533 3776 1567 3810
rect 1737 3776 1771 3810
rect 1533 3708 1567 3742
rect 1737 3708 1771 3742
rect 1533 3640 1567 3674
rect 1737 3640 1771 3674
rect 1533 3572 1567 3606
rect 1737 3572 1771 3606
rect 1533 3504 1567 3538
rect 1737 3504 1771 3538
rect 1533 3436 1567 3470
rect 1737 3436 1771 3470
rect 1533 3368 1567 3402
rect 1737 3368 1771 3402
rect 1533 3300 1567 3334
rect 1737 3300 1771 3334
rect 1533 3232 1567 3266
rect 1737 3232 1771 3266
rect 1533 3164 1567 3198
rect 1737 3164 1771 3198
rect 2095 4048 2129 4082
rect 2167 4048 2201 4082
rect 2095 3980 2129 4014
rect 2167 3980 2201 4014
rect 2095 3912 2129 3946
rect 2167 3912 2201 3946
rect 2095 3844 2129 3878
rect 2167 3844 2201 3878
rect 2095 3776 2129 3810
rect 2167 3776 2201 3810
rect 2095 3708 2129 3742
rect 2167 3708 2201 3742
rect 2095 3640 2129 3674
rect 2167 3640 2201 3674
rect 2095 3572 2129 3606
rect 2167 3572 2201 3606
rect 2095 3504 2129 3538
rect 2167 3504 2201 3538
rect 2095 3436 2129 3470
rect 2167 3436 2201 3470
rect 2095 3368 2129 3402
rect 2167 3368 2201 3402
rect 2095 3300 2129 3334
rect 2167 3300 2201 3334
rect 2095 3232 2129 3266
rect 2167 3232 2201 3266
rect 2095 3164 2129 3198
rect 2167 3164 2201 3198
rect 2525 4048 2559 4082
rect 2729 4048 2763 4082
rect 2525 3980 2559 4014
rect 2729 3980 2763 4014
rect 2525 3912 2559 3946
rect 2729 3912 2763 3946
rect 2525 3844 2559 3878
rect 2729 3844 2763 3878
rect 2525 3776 2559 3810
rect 2729 3776 2763 3810
rect 2525 3708 2559 3742
rect 2729 3708 2763 3742
rect 2525 3640 2559 3674
rect 2729 3640 2763 3674
rect 2525 3572 2559 3606
rect 2729 3572 2763 3606
rect 2525 3504 2559 3538
rect 2729 3504 2763 3538
rect 2525 3436 2559 3470
rect 2729 3436 2763 3470
rect 2525 3368 2559 3402
rect 2729 3368 2763 3402
rect 2525 3300 2559 3334
rect 2729 3300 2763 3334
rect 2525 3232 2559 3266
rect 2729 3232 2763 3266
rect 2525 3164 2559 3198
rect 2729 3164 2763 3198
rect 3087 4048 3121 4082
rect 3159 4048 3193 4082
rect 3087 3980 3121 4014
rect 3159 3980 3193 4014
rect 3087 3912 3121 3946
rect 3159 3912 3193 3946
rect 3087 3844 3121 3878
rect 3159 3844 3193 3878
rect 3087 3776 3121 3810
rect 3159 3776 3193 3810
rect 3087 3708 3121 3742
rect 3159 3708 3193 3742
rect 3087 3640 3121 3674
rect 3159 3640 3193 3674
rect 3087 3572 3121 3606
rect 3159 3572 3193 3606
rect 3087 3504 3121 3538
rect 3159 3504 3193 3538
rect 3087 3436 3121 3470
rect 3159 3436 3193 3470
rect 3087 3368 3121 3402
rect 3159 3368 3193 3402
rect 3087 3300 3121 3334
rect 3159 3300 3193 3334
rect 3087 3232 3121 3266
rect 3159 3232 3193 3266
rect 3087 3164 3121 3198
rect 3159 3164 3193 3198
rect 3517 4048 3551 4082
rect 3721 4048 3755 4082
rect 3517 3980 3551 4014
rect 3721 3980 3755 4014
rect 3517 3912 3551 3946
rect 3721 3912 3755 3946
rect 3517 3844 3551 3878
rect 3721 3844 3755 3878
rect 3517 3776 3551 3810
rect 3721 3776 3755 3810
rect 3517 3708 3551 3742
rect 3721 3708 3755 3742
rect 3517 3640 3551 3674
rect 3721 3640 3755 3674
rect 3517 3572 3551 3606
rect 3721 3572 3755 3606
rect 3517 3504 3551 3538
rect 3721 3504 3755 3538
rect 3517 3436 3551 3470
rect 3721 3436 3755 3470
rect 3517 3368 3551 3402
rect 3721 3368 3755 3402
rect 3517 3300 3551 3334
rect 3721 3300 3755 3334
rect 3517 3232 3551 3266
rect 3721 3232 3755 3266
rect 3517 3164 3551 3198
rect 3721 3164 3755 3198
rect 4079 4048 4113 4082
rect 4151 4048 4185 4082
rect 4079 3980 4113 4014
rect 4151 3980 4185 4014
rect 4079 3912 4113 3946
rect 4151 3912 4185 3946
rect 4079 3844 4113 3878
rect 4151 3844 4185 3878
rect 4079 3776 4113 3810
rect 4151 3776 4185 3810
rect 4079 3708 4113 3742
rect 4151 3708 4185 3742
rect 4079 3640 4113 3674
rect 4151 3640 4185 3674
rect 4079 3572 4113 3606
rect 4151 3572 4185 3606
rect 4079 3504 4113 3538
rect 4151 3504 4185 3538
rect 4079 3436 4113 3470
rect 4151 3436 4185 3470
rect 4079 3368 4113 3402
rect 4151 3368 4185 3402
rect 4079 3300 4113 3334
rect 4151 3300 4185 3334
rect 4079 3232 4113 3266
rect 4151 3232 4185 3266
rect 4079 3164 4113 3198
rect 4151 3164 4185 3198
rect 4509 4048 4543 4082
rect 4713 4048 4747 4082
rect 4509 3980 4543 4014
rect 4713 3980 4747 4014
rect 4509 3912 4543 3946
rect 4713 3912 4747 3946
rect 4509 3844 4543 3878
rect 4713 3844 4747 3878
rect 4509 3776 4543 3810
rect 4713 3776 4747 3810
rect 4509 3708 4543 3742
rect 4713 3708 4747 3742
rect 4509 3640 4543 3674
rect 4713 3640 4747 3674
rect 4509 3572 4543 3606
rect 4713 3572 4747 3606
rect 4509 3504 4543 3538
rect 4713 3504 4747 3538
rect 4509 3436 4543 3470
rect 4713 3436 4747 3470
rect 4509 3368 4543 3402
rect 4713 3368 4747 3402
rect 4509 3300 4543 3334
rect 4713 3300 4747 3334
rect 4509 3232 4543 3266
rect 4713 3232 4747 3266
rect 4509 3164 4543 3198
rect 4713 3164 4747 3198
rect 5071 4048 5105 4082
rect 5143 4048 5177 4082
rect 5071 3980 5105 4014
rect 5143 3980 5177 4014
rect 5071 3912 5105 3946
rect 5143 3912 5177 3946
rect 5071 3844 5105 3878
rect 5143 3844 5177 3878
rect 5071 3776 5105 3810
rect 5143 3776 5177 3810
rect 5071 3708 5105 3742
rect 5143 3708 5177 3742
rect 5071 3640 5105 3674
rect 5143 3640 5177 3674
rect 5071 3572 5105 3606
rect 5143 3572 5177 3606
rect 5071 3504 5105 3538
rect 5143 3504 5177 3538
rect 5071 3436 5105 3470
rect 5143 3436 5177 3470
rect 5071 3368 5105 3402
rect 5143 3368 5177 3402
rect 5071 3300 5105 3334
rect 5143 3300 5177 3334
rect 5071 3232 5105 3266
rect 5143 3232 5177 3266
rect 5071 3164 5105 3198
rect 5143 3164 5177 3198
rect 5501 4048 5535 4082
rect 5705 4048 5739 4082
rect 5501 3980 5535 4014
rect 5705 3980 5739 4014
rect 5501 3912 5535 3946
rect 5705 3912 5739 3946
rect 5501 3844 5535 3878
rect 5705 3844 5739 3878
rect 5501 3776 5535 3810
rect 5705 3776 5739 3810
rect 5501 3708 5535 3742
rect 5705 3708 5739 3742
rect 5501 3640 5535 3674
rect 5705 3640 5739 3674
rect 5501 3572 5535 3606
rect 5705 3572 5739 3606
rect 5501 3504 5535 3538
rect 5705 3504 5739 3538
rect 5501 3436 5535 3470
rect 5705 3436 5739 3470
rect 5501 3368 5535 3402
rect 5705 3368 5739 3402
rect 5501 3300 5535 3334
rect 5705 3300 5739 3334
rect 5501 3232 5535 3266
rect 5705 3232 5739 3266
rect 5501 3164 5535 3198
rect 5705 3164 5739 3198
rect 6063 4048 6097 4082
rect 6135 4048 6169 4082
rect 6063 3980 6097 4014
rect 6135 3980 6169 4014
rect 6063 3912 6097 3946
rect 6135 3912 6169 3946
rect 6063 3844 6097 3878
rect 6135 3844 6169 3878
rect 6063 3776 6097 3810
rect 6135 3776 6169 3810
rect 6063 3708 6097 3742
rect 6135 3708 6169 3742
rect 6063 3640 6097 3674
rect 6135 3640 6169 3674
rect 6063 3572 6097 3606
rect 6135 3572 6169 3606
rect 6063 3504 6097 3538
rect 6135 3504 6169 3538
rect 6063 3436 6097 3470
rect 6135 3436 6169 3470
rect 6063 3368 6097 3402
rect 6135 3368 6169 3402
rect 6063 3300 6097 3334
rect 6135 3300 6169 3334
rect 6063 3232 6097 3266
rect 6135 3232 6169 3266
rect 6063 3164 6097 3198
rect 6135 3164 6169 3198
rect 6493 4048 6527 4082
rect 6697 4048 6731 4082
rect 6493 3980 6527 4014
rect 6697 3980 6731 4014
rect 6493 3912 6527 3946
rect 6697 3912 6731 3946
rect 6493 3844 6527 3878
rect 6697 3844 6731 3878
rect 6493 3776 6527 3810
rect 6697 3776 6731 3810
rect 6493 3708 6527 3742
rect 6697 3708 6731 3742
rect 6493 3640 6527 3674
rect 6697 3640 6731 3674
rect 6493 3572 6527 3606
rect 6697 3572 6731 3606
rect 6493 3504 6527 3538
rect 6697 3504 6731 3538
rect 6493 3436 6527 3470
rect 6697 3436 6731 3470
rect 6493 3368 6527 3402
rect 6697 3368 6731 3402
rect 6493 3300 6527 3334
rect 6697 3300 6731 3334
rect 6493 3232 6527 3266
rect 6697 3232 6731 3266
rect 6493 3164 6527 3198
rect 6697 3164 6731 3198
rect 7055 4048 7089 4082
rect 7127 4048 7161 4082
rect 7055 3980 7089 4014
rect 7127 3980 7161 4014
rect 7055 3912 7089 3946
rect 7127 3912 7161 3946
rect 7055 3844 7089 3878
rect 7127 3844 7161 3878
rect 7055 3776 7089 3810
rect 7127 3776 7161 3810
rect 7055 3708 7089 3742
rect 7127 3708 7161 3742
rect 7055 3640 7089 3674
rect 7127 3640 7161 3674
rect 7055 3572 7089 3606
rect 7127 3572 7161 3606
rect 7055 3504 7089 3538
rect 7127 3504 7161 3538
rect 7055 3436 7089 3470
rect 7127 3436 7161 3470
rect 7055 3368 7089 3402
rect 7127 3368 7161 3402
rect 7055 3300 7089 3334
rect 7127 3300 7161 3334
rect 7055 3232 7089 3266
rect 7127 3232 7161 3266
rect 7055 3164 7089 3198
rect 7127 3164 7161 3198
rect 7485 4048 7519 4082
rect 7689 4048 7723 4082
rect 7485 3980 7519 4014
rect 7689 3980 7723 4014
rect 7485 3912 7519 3946
rect 7689 3912 7723 3946
rect 7485 3844 7519 3878
rect 7689 3844 7723 3878
rect 7485 3776 7519 3810
rect 7689 3776 7723 3810
rect 7485 3708 7519 3742
rect 7689 3708 7723 3742
rect 7485 3640 7519 3674
rect 7689 3640 7723 3674
rect 7485 3572 7519 3606
rect 7689 3572 7723 3606
rect 7485 3504 7519 3538
rect 7689 3504 7723 3538
rect 7485 3436 7519 3470
rect 7689 3436 7723 3470
rect 7485 3368 7519 3402
rect 7689 3368 7723 3402
rect 7485 3300 7519 3334
rect 7689 3300 7723 3334
rect 7485 3232 7519 3266
rect 7689 3232 7723 3266
rect 7485 3164 7519 3198
rect 7689 3164 7723 3198
rect 8047 4048 8081 4082
rect 8119 4048 8153 4082
rect 8047 3980 8081 4014
rect 8119 3980 8153 4014
rect 8047 3912 8081 3946
rect 8119 3912 8153 3946
rect 8047 3844 8081 3878
rect 8119 3844 8153 3878
rect 8047 3776 8081 3810
rect 8119 3776 8153 3810
rect 8047 3708 8081 3742
rect 8119 3708 8153 3742
rect 8047 3640 8081 3674
rect 8119 3640 8153 3674
rect 8047 3572 8081 3606
rect 8119 3572 8153 3606
rect 8047 3504 8081 3538
rect 8119 3504 8153 3538
rect 8047 3436 8081 3470
rect 8119 3436 8153 3470
rect 8047 3368 8081 3402
rect 8119 3368 8153 3402
rect 8047 3300 8081 3334
rect 8119 3300 8153 3334
rect 8047 3232 8081 3266
rect 8119 3232 8153 3266
rect 8047 3164 8081 3198
rect 8119 3164 8153 3198
rect 8477 4048 8511 4082
rect 8681 4048 8715 4082
rect 8477 3980 8511 4014
rect 8681 3980 8715 4014
rect 8477 3912 8511 3946
rect 8681 3912 8715 3946
rect 8477 3844 8511 3878
rect 8681 3844 8715 3878
rect 8477 3776 8511 3810
rect 8681 3776 8715 3810
rect 8477 3708 8511 3742
rect 8681 3708 8715 3742
rect 8477 3640 8511 3674
rect 8681 3640 8715 3674
rect 8477 3572 8511 3606
rect 8681 3572 8715 3606
rect 8477 3504 8511 3538
rect 8681 3504 8715 3538
rect 8477 3436 8511 3470
rect 8681 3436 8715 3470
rect 8477 3368 8511 3402
rect 8681 3368 8715 3402
rect 8477 3300 8511 3334
rect 8681 3300 8715 3334
rect 8477 3232 8511 3266
rect 8681 3232 8715 3266
rect 8477 3164 8511 3198
rect 8681 3164 8715 3198
rect 9039 4048 9073 4082
rect 9111 4048 9145 4082
rect 9039 3980 9073 4014
rect 9111 3980 9145 4014
rect 9039 3912 9073 3946
rect 9111 3912 9145 3946
rect 9039 3844 9073 3878
rect 9111 3844 9145 3878
rect 9039 3776 9073 3810
rect 9111 3776 9145 3810
rect 9039 3708 9073 3742
rect 9111 3708 9145 3742
rect 9039 3640 9073 3674
rect 9111 3640 9145 3674
rect 9039 3572 9073 3606
rect 9111 3572 9145 3606
rect 9039 3504 9073 3538
rect 9111 3504 9145 3538
rect 9039 3436 9073 3470
rect 9111 3436 9145 3470
rect 9039 3368 9073 3402
rect 9111 3368 9145 3402
rect 9039 3300 9073 3334
rect 9111 3300 9145 3334
rect 9039 3232 9073 3266
rect 9111 3232 9145 3266
rect 9039 3164 9073 3198
rect 9111 3164 9145 3198
rect 9469 4048 9503 4082
rect 9673 4048 9707 4082
rect 9469 3980 9503 4014
rect 9673 3980 9707 4014
rect 9469 3912 9503 3946
rect 9673 3912 9707 3946
rect 9469 3844 9503 3878
rect 9673 3844 9707 3878
rect 9469 3776 9503 3810
rect 9673 3776 9707 3810
rect 9469 3708 9503 3742
rect 9673 3708 9707 3742
rect 9469 3640 9503 3674
rect 9673 3640 9707 3674
rect 9469 3572 9503 3606
rect 9673 3572 9707 3606
rect 9469 3504 9503 3538
rect 9673 3504 9707 3538
rect 9469 3436 9503 3470
rect 9673 3436 9707 3470
rect 9469 3368 9503 3402
rect 9673 3368 9707 3402
rect 9469 3300 9503 3334
rect 9673 3300 9707 3334
rect 9469 3232 9503 3266
rect 9673 3232 9707 3266
rect 9469 3164 9503 3198
rect 9673 3164 9707 3198
rect 10031 4048 10065 4082
rect 10103 4048 10137 4082
rect 10031 3980 10065 4014
rect 10103 3980 10137 4014
rect 10031 3912 10065 3946
rect 10103 3912 10137 3946
rect 10031 3844 10065 3878
rect 10103 3844 10137 3878
rect 10031 3776 10065 3810
rect 10103 3776 10137 3810
rect 10031 3708 10065 3742
rect 10103 3708 10137 3742
rect 10031 3640 10065 3674
rect 10103 3640 10137 3674
rect 10031 3572 10065 3606
rect 10103 3572 10137 3606
rect 10031 3504 10065 3538
rect 10103 3504 10137 3538
rect 10031 3436 10065 3470
rect 10103 3436 10137 3470
rect 10031 3368 10065 3402
rect 10103 3368 10137 3402
rect 10031 3300 10065 3334
rect 10103 3300 10137 3334
rect 10031 3232 10065 3266
rect 10103 3232 10137 3266
rect 10031 3164 10065 3198
rect 10103 3164 10137 3198
rect 10461 4048 10495 4082
rect 10665 4048 10699 4082
rect 10461 3980 10495 4014
rect 10665 3980 10699 4014
rect 10461 3912 10495 3946
rect 10665 3912 10699 3946
rect 10461 3844 10495 3878
rect 10665 3844 10699 3878
rect 10461 3776 10495 3810
rect 10665 3776 10699 3810
rect 10461 3708 10495 3742
rect 10665 3708 10699 3742
rect 10461 3640 10495 3674
rect 10665 3640 10699 3674
rect 10461 3572 10495 3606
rect 10665 3572 10699 3606
rect 10461 3504 10495 3538
rect 10665 3504 10699 3538
rect 10461 3436 10495 3470
rect 10665 3436 10699 3470
rect 10461 3368 10495 3402
rect 10665 3368 10699 3402
rect 10461 3300 10495 3334
rect 10665 3300 10699 3334
rect 10461 3232 10495 3266
rect 10665 3232 10699 3266
rect 10461 3164 10495 3198
rect 10665 3164 10699 3198
rect 11023 4048 11057 4082
rect 11095 4048 11129 4082
rect 11023 3980 11057 4014
rect 11095 3980 11129 4014
rect 11023 3912 11057 3946
rect 11095 3912 11129 3946
rect 11023 3844 11057 3878
rect 11095 3844 11129 3878
rect 11023 3776 11057 3810
rect 11095 3776 11129 3810
rect 11023 3708 11057 3742
rect 11095 3708 11129 3742
rect 11023 3640 11057 3674
rect 11095 3640 11129 3674
rect 11023 3572 11057 3606
rect 11095 3572 11129 3606
rect 11023 3504 11057 3538
rect 11095 3504 11129 3538
rect 11023 3436 11057 3470
rect 11095 3436 11129 3470
rect 11023 3368 11057 3402
rect 11095 3368 11129 3402
rect 11023 3300 11057 3334
rect 11095 3300 11129 3334
rect 11023 3232 11057 3266
rect 11095 3232 11129 3266
rect 11023 3164 11057 3198
rect 11095 3164 11129 3198
rect 11453 4048 11487 4082
rect 11657 4048 11691 4082
rect 11453 3980 11487 4014
rect 11657 3980 11691 4014
rect 11453 3912 11487 3946
rect 11657 3912 11691 3946
rect 11453 3844 11487 3878
rect 11657 3844 11691 3878
rect 11453 3776 11487 3810
rect 11657 3776 11691 3810
rect 11453 3708 11487 3742
rect 11657 3708 11691 3742
rect 11453 3640 11487 3674
rect 11657 3640 11691 3674
rect 11453 3572 11487 3606
rect 11657 3572 11691 3606
rect 11453 3504 11487 3538
rect 11657 3504 11691 3538
rect 11453 3436 11487 3470
rect 11657 3436 11691 3470
rect 11453 3368 11487 3402
rect 11657 3368 11691 3402
rect 11453 3300 11487 3334
rect 11657 3300 11691 3334
rect 11453 3232 11487 3266
rect 11657 3232 11691 3266
rect 11453 3164 11487 3198
rect 11657 3164 11691 3198
rect 12015 4048 12049 4082
rect 12087 4048 12121 4082
rect 12015 3980 12049 4014
rect 12087 3980 12121 4014
rect 12015 3912 12049 3946
rect 12087 3912 12121 3946
rect 12015 3844 12049 3878
rect 12087 3844 12121 3878
rect 12015 3776 12049 3810
rect 12087 3776 12121 3810
rect 12015 3708 12049 3742
rect 12087 3708 12121 3742
rect 12015 3640 12049 3674
rect 12087 3640 12121 3674
rect 12015 3572 12049 3606
rect 12087 3572 12121 3606
rect 12015 3504 12049 3538
rect 12087 3504 12121 3538
rect 12015 3436 12049 3470
rect 12087 3436 12121 3470
rect 12015 3368 12049 3402
rect 12087 3368 12121 3402
rect 12015 3300 12049 3334
rect 12087 3300 12121 3334
rect 12015 3232 12049 3266
rect 12087 3232 12121 3266
rect 12015 3164 12049 3198
rect 12087 3164 12121 3198
rect 12445 4048 12479 4082
rect 12649 4048 12683 4082
rect 12445 3980 12479 4014
rect 12649 3980 12683 4014
rect 12445 3912 12479 3946
rect 12649 3912 12683 3946
rect 12445 3844 12479 3878
rect 12649 3844 12683 3878
rect 12445 3776 12479 3810
rect 12649 3776 12683 3810
rect 12445 3708 12479 3742
rect 12649 3708 12683 3742
rect 12445 3640 12479 3674
rect 12649 3640 12683 3674
rect 12445 3572 12479 3606
rect 12649 3572 12683 3606
rect 12445 3504 12479 3538
rect 12649 3504 12683 3538
rect 12445 3436 12479 3470
rect 12649 3436 12683 3470
rect 12445 3368 12479 3402
rect 12649 3368 12683 3402
rect 12445 3300 12479 3334
rect 12649 3300 12683 3334
rect 12445 3232 12479 3266
rect 12649 3232 12683 3266
rect 12445 3164 12479 3198
rect 12649 3164 12683 3198
rect 13007 4048 13041 4082
rect 13079 4048 13113 4082
rect 13007 3980 13041 4014
rect 13079 3980 13113 4014
rect 13007 3912 13041 3946
rect 13079 3912 13113 3946
rect 13007 3844 13041 3878
rect 13079 3844 13113 3878
rect 13007 3776 13041 3810
rect 13079 3776 13113 3810
rect 13007 3708 13041 3742
rect 13079 3708 13113 3742
rect 13007 3640 13041 3674
rect 13079 3640 13113 3674
rect 13007 3572 13041 3606
rect 13079 3572 13113 3606
rect 13007 3504 13041 3538
rect 13079 3504 13113 3538
rect 13007 3436 13041 3470
rect 13079 3436 13113 3470
rect 13007 3368 13041 3402
rect 13079 3368 13113 3402
rect 13007 3300 13041 3334
rect 13079 3300 13113 3334
rect 13007 3232 13041 3266
rect 13079 3232 13113 3266
rect 13007 3164 13041 3198
rect 13079 3164 13113 3198
rect 13437 4048 13471 4082
rect 13641 4048 13675 4082
rect 13437 3980 13471 4014
rect 13641 3980 13675 4014
rect 13437 3912 13471 3946
rect 13641 3912 13675 3946
rect 13437 3844 13471 3878
rect 13641 3844 13675 3878
rect 13437 3776 13471 3810
rect 13641 3776 13675 3810
rect 13437 3708 13471 3742
rect 13641 3708 13675 3742
rect 13437 3640 13471 3674
rect 13641 3640 13675 3674
rect 13437 3572 13471 3606
rect 13641 3572 13675 3606
rect 13437 3504 13471 3538
rect 13641 3504 13675 3538
rect 13437 3436 13471 3470
rect 13641 3436 13675 3470
rect 13437 3368 13471 3402
rect 13641 3368 13675 3402
rect 13437 3300 13471 3334
rect 13641 3300 13675 3334
rect 13437 3232 13471 3266
rect 13641 3232 13675 3266
rect 13437 3164 13471 3198
rect 13641 3164 13675 3198
rect 13999 4048 14033 4082
rect 13999 3980 14033 4014
rect 13999 3912 14033 3946
rect 13999 3844 14033 3878
rect 13999 3776 14033 3810
rect 13999 3708 14033 3742
rect 13999 3640 14033 3674
rect 13999 3572 14033 3606
rect 13999 3504 14033 3538
rect 13999 3436 14033 3470
rect 13999 3368 14033 3402
rect 13999 3300 14033 3334
rect 13999 3232 14033 3266
rect 13999 3164 14033 3198
rect 14356 4048 14390 4082
rect 14356 3980 14390 4014
rect 14356 3912 14390 3946
rect 14356 3844 14390 3878
rect 14356 3776 14390 3810
rect 14356 3708 14390 3742
rect 14356 3640 14390 3674
rect 14356 3572 14390 3606
rect 14356 3504 14390 3538
rect 14356 3436 14390 3470
rect 14356 3368 14390 3402
rect 14356 3300 14390 3334
rect 14356 3232 14390 3266
rect 14356 3164 14390 3198
rect 745 2448 779 2482
rect 745 2380 779 2414
rect 745 2312 779 2346
rect 745 2244 779 2278
rect 745 2176 779 2210
rect 745 2108 779 2142
rect 745 2040 779 2074
rect 745 1972 779 2006
rect 745 1904 779 1938
rect 745 1836 779 1870
rect 745 1768 779 1802
rect 745 1700 779 1734
rect 745 1632 779 1666
rect 745 1564 779 1598
rect 1103 2448 1137 2482
rect 1175 2448 1209 2482
rect 1103 2380 1137 2414
rect 1175 2380 1209 2414
rect 1103 2312 1137 2346
rect 1175 2312 1209 2346
rect 1103 2244 1137 2278
rect 1175 2244 1209 2278
rect 1103 2176 1137 2210
rect 1175 2176 1209 2210
rect 1103 2108 1137 2142
rect 1175 2108 1209 2142
rect 1103 2040 1137 2074
rect 1175 2040 1209 2074
rect 1103 1972 1137 2006
rect 1175 1972 1209 2006
rect 1103 1904 1137 1938
rect 1175 1904 1209 1938
rect 1103 1836 1137 1870
rect 1175 1836 1209 1870
rect 1103 1768 1137 1802
rect 1175 1768 1209 1802
rect 1103 1700 1137 1734
rect 1175 1700 1209 1734
rect 1103 1632 1137 1666
rect 1175 1632 1209 1666
rect 1103 1564 1137 1598
rect 1175 1564 1209 1598
rect 1533 2506 1567 2540
rect 1737 2506 1771 2540
rect 1533 2438 1567 2472
rect 1737 2438 1771 2472
rect 1533 2370 1567 2404
rect 1737 2370 1771 2404
rect 1533 2302 1567 2336
rect 1737 2302 1771 2336
rect 1533 2234 1567 2268
rect 1737 2234 1771 2268
rect 1533 2166 1567 2200
rect 1737 2166 1771 2200
rect 1533 2098 1567 2132
rect 1737 2098 1771 2132
rect 1533 2030 1567 2064
rect 1737 2030 1771 2064
rect 1533 1962 1567 1996
rect 1737 1962 1771 1996
rect 1533 1894 1567 1928
rect 1737 1894 1771 1928
rect 1533 1826 1567 1860
rect 1737 1826 1771 1860
rect 1533 1758 1567 1792
rect 1737 1758 1771 1792
rect 1533 1690 1567 1724
rect 1737 1690 1771 1724
rect 1533 1622 1567 1656
rect 1737 1622 1771 1656
rect 2095 2448 2129 2482
rect 2167 2448 2201 2482
rect 2095 2380 2129 2414
rect 2167 2380 2201 2414
rect 2095 2312 2129 2346
rect 2167 2312 2201 2346
rect 2095 2244 2129 2278
rect 2167 2244 2201 2278
rect 2095 2176 2129 2210
rect 2167 2176 2201 2210
rect 2095 2108 2129 2142
rect 2167 2108 2201 2142
rect 2095 2040 2129 2074
rect 2167 2040 2201 2074
rect 2095 1972 2129 2006
rect 2167 1972 2201 2006
rect 2095 1904 2129 1938
rect 2167 1904 2201 1938
rect 2095 1836 2129 1870
rect 2167 1836 2201 1870
rect 2095 1768 2129 1802
rect 2167 1768 2201 1802
rect 2095 1700 2129 1734
rect 2167 1700 2201 1734
rect 2095 1632 2129 1666
rect 2167 1632 2201 1666
rect 2095 1564 2129 1598
rect 2167 1564 2201 1598
rect 2525 2506 2559 2540
rect 2729 2506 2763 2540
rect 2525 2438 2559 2472
rect 2729 2438 2763 2472
rect 2525 2370 2559 2404
rect 2729 2370 2763 2404
rect 2525 2302 2559 2336
rect 2729 2302 2763 2336
rect 2525 2234 2559 2268
rect 2729 2234 2763 2268
rect 2525 2166 2559 2200
rect 2729 2166 2763 2200
rect 2525 2098 2559 2132
rect 2729 2098 2763 2132
rect 2525 2030 2559 2064
rect 2729 2030 2763 2064
rect 2525 1962 2559 1996
rect 2729 1962 2763 1996
rect 2525 1894 2559 1928
rect 2729 1894 2763 1928
rect 2525 1826 2559 1860
rect 2729 1826 2763 1860
rect 2525 1758 2559 1792
rect 2729 1758 2763 1792
rect 2525 1690 2559 1724
rect 2729 1690 2763 1724
rect 2525 1622 2559 1656
rect 2729 1622 2763 1656
rect 3087 2448 3121 2482
rect 3159 2448 3193 2482
rect 3087 2380 3121 2414
rect 3159 2380 3193 2414
rect 3087 2312 3121 2346
rect 3159 2312 3193 2346
rect 3087 2244 3121 2278
rect 3159 2244 3193 2278
rect 3087 2176 3121 2210
rect 3159 2176 3193 2210
rect 3087 2108 3121 2142
rect 3159 2108 3193 2142
rect 3087 2040 3121 2074
rect 3159 2040 3193 2074
rect 3087 1972 3121 2006
rect 3159 1972 3193 2006
rect 3087 1904 3121 1938
rect 3159 1904 3193 1938
rect 3087 1836 3121 1870
rect 3159 1836 3193 1870
rect 3087 1768 3121 1802
rect 3159 1768 3193 1802
rect 3087 1700 3121 1734
rect 3159 1700 3193 1734
rect 3087 1632 3121 1666
rect 3159 1632 3193 1666
rect 3087 1564 3121 1598
rect 3159 1564 3193 1598
rect 3517 2506 3551 2540
rect 3721 2506 3755 2540
rect 3517 2438 3551 2472
rect 3721 2438 3755 2472
rect 3517 2370 3551 2404
rect 3721 2370 3755 2404
rect 3517 2302 3551 2336
rect 3721 2302 3755 2336
rect 3517 2234 3551 2268
rect 3721 2234 3755 2268
rect 3517 2166 3551 2200
rect 3721 2166 3755 2200
rect 3517 2098 3551 2132
rect 3721 2098 3755 2132
rect 3517 2030 3551 2064
rect 3721 2030 3755 2064
rect 3517 1962 3551 1996
rect 3721 1962 3755 1996
rect 3517 1894 3551 1928
rect 3721 1894 3755 1928
rect 3517 1826 3551 1860
rect 3721 1826 3755 1860
rect 3517 1758 3551 1792
rect 3721 1758 3755 1792
rect 3517 1690 3551 1724
rect 3721 1690 3755 1724
rect 3517 1622 3551 1656
rect 3721 1622 3755 1656
rect 4079 2448 4113 2482
rect 4151 2448 4185 2482
rect 4079 2380 4113 2414
rect 4151 2380 4185 2414
rect 4079 2312 4113 2346
rect 4151 2312 4185 2346
rect 4079 2244 4113 2278
rect 4151 2244 4185 2278
rect 4079 2176 4113 2210
rect 4151 2176 4185 2210
rect 4079 2108 4113 2142
rect 4151 2108 4185 2142
rect 4079 2040 4113 2074
rect 4151 2040 4185 2074
rect 4079 1972 4113 2006
rect 4151 1972 4185 2006
rect 4079 1904 4113 1938
rect 4151 1904 4185 1938
rect 4079 1836 4113 1870
rect 4151 1836 4185 1870
rect 4079 1768 4113 1802
rect 4151 1768 4185 1802
rect 4079 1700 4113 1734
rect 4151 1700 4185 1734
rect 4079 1632 4113 1666
rect 4151 1632 4185 1666
rect 4079 1564 4113 1598
rect 4151 1564 4185 1598
rect 4509 2506 4543 2540
rect 4713 2506 4747 2540
rect 4509 2438 4543 2472
rect 4713 2438 4747 2472
rect 4509 2370 4543 2404
rect 4713 2370 4747 2404
rect 4509 2302 4543 2336
rect 4713 2302 4747 2336
rect 4509 2234 4543 2268
rect 4713 2234 4747 2268
rect 4509 2166 4543 2200
rect 4713 2166 4747 2200
rect 4509 2098 4543 2132
rect 4713 2098 4747 2132
rect 4509 2030 4543 2064
rect 4713 2030 4747 2064
rect 4509 1962 4543 1996
rect 4713 1962 4747 1996
rect 4509 1894 4543 1928
rect 4713 1894 4747 1928
rect 4509 1826 4543 1860
rect 4713 1826 4747 1860
rect 4509 1758 4543 1792
rect 4713 1758 4747 1792
rect 4509 1690 4543 1724
rect 4713 1690 4747 1724
rect 4509 1622 4543 1656
rect 4713 1622 4747 1656
rect 5071 2448 5105 2482
rect 5143 2448 5177 2482
rect 5071 2380 5105 2414
rect 5143 2380 5177 2414
rect 5071 2312 5105 2346
rect 5143 2312 5177 2346
rect 5071 2244 5105 2278
rect 5143 2244 5177 2278
rect 5071 2176 5105 2210
rect 5143 2176 5177 2210
rect 5071 2108 5105 2142
rect 5143 2108 5177 2142
rect 5071 2040 5105 2074
rect 5143 2040 5177 2074
rect 5071 1972 5105 2006
rect 5143 1972 5177 2006
rect 5071 1904 5105 1938
rect 5143 1904 5177 1938
rect 5071 1836 5105 1870
rect 5143 1836 5177 1870
rect 5071 1768 5105 1802
rect 5143 1768 5177 1802
rect 5071 1700 5105 1734
rect 5143 1700 5177 1734
rect 5071 1632 5105 1666
rect 5143 1632 5177 1666
rect 5071 1564 5105 1598
rect 5143 1564 5177 1598
rect 5501 2506 5535 2540
rect 5705 2506 5739 2540
rect 5501 2438 5535 2472
rect 5705 2438 5739 2472
rect 5501 2370 5535 2404
rect 5705 2370 5739 2404
rect 5501 2302 5535 2336
rect 5705 2302 5739 2336
rect 5501 2234 5535 2268
rect 5705 2234 5739 2268
rect 5501 2166 5535 2200
rect 5705 2166 5739 2200
rect 5501 2098 5535 2132
rect 5705 2098 5739 2132
rect 5501 2030 5535 2064
rect 5705 2030 5739 2064
rect 5501 1962 5535 1996
rect 5705 1962 5739 1996
rect 5501 1894 5535 1928
rect 5705 1894 5739 1928
rect 5501 1826 5535 1860
rect 5705 1826 5739 1860
rect 5501 1758 5535 1792
rect 5705 1758 5739 1792
rect 5501 1690 5535 1724
rect 5705 1690 5739 1724
rect 5501 1622 5535 1656
rect 5705 1622 5739 1656
rect 6063 2448 6097 2482
rect 6135 2448 6169 2482
rect 6063 2380 6097 2414
rect 6135 2380 6169 2414
rect 6063 2312 6097 2346
rect 6135 2312 6169 2346
rect 6063 2244 6097 2278
rect 6135 2244 6169 2278
rect 6063 2176 6097 2210
rect 6135 2176 6169 2210
rect 6063 2108 6097 2142
rect 6135 2108 6169 2142
rect 6063 2040 6097 2074
rect 6135 2040 6169 2074
rect 6063 1972 6097 2006
rect 6135 1972 6169 2006
rect 6063 1904 6097 1938
rect 6135 1904 6169 1938
rect 6063 1836 6097 1870
rect 6135 1836 6169 1870
rect 6063 1768 6097 1802
rect 6135 1768 6169 1802
rect 6063 1700 6097 1734
rect 6135 1700 6169 1734
rect 6063 1632 6097 1666
rect 6135 1632 6169 1666
rect 6063 1564 6097 1598
rect 6135 1564 6169 1598
rect 6493 2506 6527 2540
rect 6697 2506 6731 2540
rect 6493 2438 6527 2472
rect 6697 2438 6731 2472
rect 6493 2370 6527 2404
rect 6697 2370 6731 2404
rect 6493 2302 6527 2336
rect 6697 2302 6731 2336
rect 6493 2234 6527 2268
rect 6697 2234 6731 2268
rect 6493 2166 6527 2200
rect 6697 2166 6731 2200
rect 6493 2098 6527 2132
rect 6697 2098 6731 2132
rect 6493 2030 6527 2064
rect 6697 2030 6731 2064
rect 6493 1962 6527 1996
rect 6697 1962 6731 1996
rect 6493 1894 6527 1928
rect 6697 1894 6731 1928
rect 6493 1826 6527 1860
rect 6697 1826 6731 1860
rect 6493 1758 6527 1792
rect 6697 1758 6731 1792
rect 6493 1690 6527 1724
rect 6697 1690 6731 1724
rect 6493 1622 6527 1656
rect 6697 1622 6731 1656
rect 7055 2448 7089 2482
rect 7127 2448 7161 2482
rect 7055 2380 7089 2414
rect 7127 2380 7161 2414
rect 7055 2312 7089 2346
rect 7127 2312 7161 2346
rect 7055 2244 7089 2278
rect 7127 2244 7161 2278
rect 7055 2176 7089 2210
rect 7127 2176 7161 2210
rect 7055 2108 7089 2142
rect 7127 2108 7161 2142
rect 7055 2040 7089 2074
rect 7127 2040 7161 2074
rect 7055 1972 7089 2006
rect 7127 1972 7161 2006
rect 7055 1904 7089 1938
rect 7127 1904 7161 1938
rect 7055 1836 7089 1870
rect 7127 1836 7161 1870
rect 7055 1768 7089 1802
rect 7127 1768 7161 1802
rect 7055 1700 7089 1734
rect 7127 1700 7161 1734
rect 7055 1632 7089 1666
rect 7127 1632 7161 1666
rect 7055 1564 7089 1598
rect 7127 1564 7161 1598
rect 7485 2506 7519 2540
rect 7689 2506 7723 2540
rect 7485 2438 7519 2472
rect 7689 2438 7723 2472
rect 7485 2370 7519 2404
rect 7689 2370 7723 2404
rect 7485 2302 7519 2336
rect 7689 2302 7723 2336
rect 7485 2234 7519 2268
rect 7689 2234 7723 2268
rect 7485 2166 7519 2200
rect 7689 2166 7723 2200
rect 7485 2098 7519 2132
rect 7689 2098 7723 2132
rect 7485 2030 7519 2064
rect 7689 2030 7723 2064
rect 7485 1962 7519 1996
rect 7689 1962 7723 1996
rect 7485 1894 7519 1928
rect 7689 1894 7723 1928
rect 7485 1826 7519 1860
rect 7689 1826 7723 1860
rect 7485 1758 7519 1792
rect 7689 1758 7723 1792
rect 7485 1690 7519 1724
rect 7689 1690 7723 1724
rect 7485 1622 7519 1656
rect 7689 1622 7723 1656
rect 8047 2448 8081 2482
rect 8119 2448 8153 2482
rect 8047 2380 8081 2414
rect 8119 2380 8153 2414
rect 8047 2312 8081 2346
rect 8119 2312 8153 2346
rect 8047 2244 8081 2278
rect 8119 2244 8153 2278
rect 8047 2176 8081 2210
rect 8119 2176 8153 2210
rect 8047 2108 8081 2142
rect 8119 2108 8153 2142
rect 8047 2040 8081 2074
rect 8119 2040 8153 2074
rect 8047 1972 8081 2006
rect 8119 1972 8153 2006
rect 8047 1904 8081 1938
rect 8119 1904 8153 1938
rect 8047 1836 8081 1870
rect 8119 1836 8153 1870
rect 8047 1768 8081 1802
rect 8119 1768 8153 1802
rect 8047 1700 8081 1734
rect 8119 1700 8153 1734
rect 8047 1632 8081 1666
rect 8119 1632 8153 1666
rect 8047 1564 8081 1598
rect 8119 1564 8153 1598
rect 8477 2506 8511 2540
rect 8681 2506 8715 2540
rect 8477 2438 8511 2472
rect 8681 2438 8715 2472
rect 8477 2370 8511 2404
rect 8681 2370 8715 2404
rect 8477 2302 8511 2336
rect 8681 2302 8715 2336
rect 8477 2234 8511 2268
rect 8681 2234 8715 2268
rect 8477 2166 8511 2200
rect 8681 2166 8715 2200
rect 8477 2098 8511 2132
rect 8681 2098 8715 2132
rect 8477 2030 8511 2064
rect 8681 2030 8715 2064
rect 8477 1962 8511 1996
rect 8681 1962 8715 1996
rect 8477 1894 8511 1928
rect 8681 1894 8715 1928
rect 8477 1826 8511 1860
rect 8681 1826 8715 1860
rect 8477 1758 8511 1792
rect 8681 1758 8715 1792
rect 8477 1690 8511 1724
rect 8681 1690 8715 1724
rect 8477 1622 8511 1656
rect 8681 1622 8715 1656
rect 9039 2448 9073 2482
rect 9111 2448 9145 2482
rect 9039 2380 9073 2414
rect 9111 2380 9145 2414
rect 9039 2312 9073 2346
rect 9111 2312 9145 2346
rect 9039 2244 9073 2278
rect 9111 2244 9145 2278
rect 9039 2176 9073 2210
rect 9111 2176 9145 2210
rect 9039 2108 9073 2142
rect 9111 2108 9145 2142
rect 9039 2040 9073 2074
rect 9111 2040 9145 2074
rect 9039 1972 9073 2006
rect 9111 1972 9145 2006
rect 9039 1904 9073 1938
rect 9111 1904 9145 1938
rect 9039 1836 9073 1870
rect 9111 1836 9145 1870
rect 9039 1768 9073 1802
rect 9111 1768 9145 1802
rect 9039 1700 9073 1734
rect 9111 1700 9145 1734
rect 9039 1632 9073 1666
rect 9111 1632 9145 1666
rect 9039 1564 9073 1598
rect 9111 1564 9145 1598
rect 9469 2506 9503 2540
rect 9673 2506 9707 2540
rect 9469 2438 9503 2472
rect 9673 2438 9707 2472
rect 9469 2370 9503 2404
rect 9673 2370 9707 2404
rect 9469 2302 9503 2336
rect 9673 2302 9707 2336
rect 9469 2234 9503 2268
rect 9673 2234 9707 2268
rect 9469 2166 9503 2200
rect 9673 2166 9707 2200
rect 9469 2098 9503 2132
rect 9673 2098 9707 2132
rect 9469 2030 9503 2064
rect 9673 2030 9707 2064
rect 9469 1962 9503 1996
rect 9673 1962 9707 1996
rect 9469 1894 9503 1928
rect 9673 1894 9707 1928
rect 9469 1826 9503 1860
rect 9673 1826 9707 1860
rect 9469 1758 9503 1792
rect 9673 1758 9707 1792
rect 9469 1690 9503 1724
rect 9673 1690 9707 1724
rect 9469 1622 9503 1656
rect 9673 1622 9707 1656
rect 10031 2448 10065 2482
rect 10103 2448 10137 2482
rect 10031 2380 10065 2414
rect 10103 2380 10137 2414
rect 10031 2312 10065 2346
rect 10103 2312 10137 2346
rect 10031 2244 10065 2278
rect 10103 2244 10137 2278
rect 10031 2176 10065 2210
rect 10103 2176 10137 2210
rect 10031 2108 10065 2142
rect 10103 2108 10137 2142
rect 10031 2040 10065 2074
rect 10103 2040 10137 2074
rect 10031 1972 10065 2006
rect 10103 1972 10137 2006
rect 10031 1904 10065 1938
rect 10103 1904 10137 1938
rect 10031 1836 10065 1870
rect 10103 1836 10137 1870
rect 10031 1768 10065 1802
rect 10103 1768 10137 1802
rect 10031 1700 10065 1734
rect 10103 1700 10137 1734
rect 10031 1632 10065 1666
rect 10103 1632 10137 1666
rect 10031 1564 10065 1598
rect 10103 1564 10137 1598
rect 10461 2506 10495 2540
rect 10665 2506 10699 2540
rect 10461 2438 10495 2472
rect 10665 2438 10699 2472
rect 10461 2370 10495 2404
rect 10665 2370 10699 2404
rect 10461 2302 10495 2336
rect 10665 2302 10699 2336
rect 10461 2234 10495 2268
rect 10665 2234 10699 2268
rect 10461 2166 10495 2200
rect 10665 2166 10699 2200
rect 10461 2098 10495 2132
rect 10665 2098 10699 2132
rect 10461 2030 10495 2064
rect 10665 2030 10699 2064
rect 10461 1962 10495 1996
rect 10665 1962 10699 1996
rect 10461 1894 10495 1928
rect 10665 1894 10699 1928
rect 10461 1826 10495 1860
rect 10665 1826 10699 1860
rect 10461 1758 10495 1792
rect 10665 1758 10699 1792
rect 10461 1690 10495 1724
rect 10665 1690 10699 1724
rect 10461 1622 10495 1656
rect 10665 1622 10699 1656
rect 11023 2448 11057 2482
rect 11095 2448 11129 2482
rect 11023 2380 11057 2414
rect 11095 2380 11129 2414
rect 11023 2312 11057 2346
rect 11095 2312 11129 2346
rect 11023 2244 11057 2278
rect 11095 2244 11129 2278
rect 11023 2176 11057 2210
rect 11095 2176 11129 2210
rect 11023 2108 11057 2142
rect 11095 2108 11129 2142
rect 11023 2040 11057 2074
rect 11095 2040 11129 2074
rect 11023 1972 11057 2006
rect 11095 1972 11129 2006
rect 11023 1904 11057 1938
rect 11095 1904 11129 1938
rect 11023 1836 11057 1870
rect 11095 1836 11129 1870
rect 11023 1768 11057 1802
rect 11095 1768 11129 1802
rect 11023 1700 11057 1734
rect 11095 1700 11129 1734
rect 11023 1632 11057 1666
rect 11095 1632 11129 1666
rect 11023 1564 11057 1598
rect 11095 1564 11129 1598
rect 11453 2506 11487 2540
rect 11657 2506 11691 2540
rect 11453 2438 11487 2472
rect 11657 2438 11691 2472
rect 11453 2370 11487 2404
rect 11657 2370 11691 2404
rect 11453 2302 11487 2336
rect 11657 2302 11691 2336
rect 11453 2234 11487 2268
rect 11657 2234 11691 2268
rect 11453 2166 11487 2200
rect 11657 2166 11691 2200
rect 11453 2098 11487 2132
rect 11657 2098 11691 2132
rect 11453 2030 11487 2064
rect 11657 2030 11691 2064
rect 11453 1962 11487 1996
rect 11657 1962 11691 1996
rect 11453 1894 11487 1928
rect 11657 1894 11691 1928
rect 11453 1826 11487 1860
rect 11657 1826 11691 1860
rect 11453 1758 11487 1792
rect 11657 1758 11691 1792
rect 11453 1690 11487 1724
rect 11657 1690 11691 1724
rect 11453 1622 11487 1656
rect 11657 1622 11691 1656
rect 12015 2448 12049 2482
rect 12087 2448 12121 2482
rect 12015 2380 12049 2414
rect 12087 2380 12121 2414
rect 12015 2312 12049 2346
rect 12087 2312 12121 2346
rect 12015 2244 12049 2278
rect 12087 2244 12121 2278
rect 12015 2176 12049 2210
rect 12087 2176 12121 2210
rect 12015 2108 12049 2142
rect 12087 2108 12121 2142
rect 12015 2040 12049 2074
rect 12087 2040 12121 2074
rect 12015 1972 12049 2006
rect 12087 1972 12121 2006
rect 12015 1904 12049 1938
rect 12087 1904 12121 1938
rect 12015 1836 12049 1870
rect 12087 1836 12121 1870
rect 12015 1768 12049 1802
rect 12087 1768 12121 1802
rect 12015 1700 12049 1734
rect 12087 1700 12121 1734
rect 12015 1632 12049 1666
rect 12087 1632 12121 1666
rect 12015 1564 12049 1598
rect 12087 1564 12121 1598
rect 12445 2506 12479 2540
rect 12649 2506 12683 2540
rect 12445 2438 12479 2472
rect 12649 2438 12683 2472
rect 12445 2370 12479 2404
rect 12649 2370 12683 2404
rect 12445 2302 12479 2336
rect 12649 2302 12683 2336
rect 12445 2234 12479 2268
rect 12649 2234 12683 2268
rect 12445 2166 12479 2200
rect 12649 2166 12683 2200
rect 12445 2098 12479 2132
rect 12649 2098 12683 2132
rect 12445 2030 12479 2064
rect 12649 2030 12683 2064
rect 12445 1962 12479 1996
rect 12649 1962 12683 1996
rect 12445 1894 12479 1928
rect 12649 1894 12683 1928
rect 12445 1826 12479 1860
rect 12649 1826 12683 1860
rect 12445 1758 12479 1792
rect 12649 1758 12683 1792
rect 12445 1690 12479 1724
rect 12649 1690 12683 1724
rect 12445 1622 12479 1656
rect 12649 1622 12683 1656
rect 13007 2448 13041 2482
rect 13079 2448 13113 2482
rect 13007 2380 13041 2414
rect 13079 2380 13113 2414
rect 13007 2312 13041 2346
rect 13079 2312 13113 2346
rect 13007 2244 13041 2278
rect 13079 2244 13113 2278
rect 13007 2176 13041 2210
rect 13079 2176 13113 2210
rect 13007 2108 13041 2142
rect 13079 2108 13113 2142
rect 13007 2040 13041 2074
rect 13079 2040 13113 2074
rect 13007 1972 13041 2006
rect 13079 1972 13113 2006
rect 13007 1904 13041 1938
rect 13079 1904 13113 1938
rect 13007 1836 13041 1870
rect 13079 1836 13113 1870
rect 13007 1768 13041 1802
rect 13079 1768 13113 1802
rect 13007 1700 13041 1734
rect 13079 1700 13113 1734
rect 13007 1632 13041 1666
rect 13079 1632 13113 1666
rect 13007 1564 13041 1598
rect 13079 1564 13113 1598
rect 13437 2506 13471 2540
rect 13641 2506 13675 2540
rect 13437 2438 13471 2472
rect 13641 2438 13675 2472
rect 13437 2370 13471 2404
rect 13641 2370 13675 2404
rect 13437 2302 13471 2336
rect 13641 2302 13675 2336
rect 13437 2234 13471 2268
rect 13641 2234 13675 2268
rect 13437 2166 13471 2200
rect 13641 2166 13675 2200
rect 13437 2098 13471 2132
rect 13641 2098 13675 2132
rect 13437 2030 13471 2064
rect 13641 2030 13675 2064
rect 13437 1962 13471 1996
rect 13641 1962 13675 1996
rect 13437 1894 13471 1928
rect 13641 1894 13675 1928
rect 13437 1826 13471 1860
rect 13641 1826 13675 1860
rect 13437 1758 13471 1792
rect 13641 1758 13675 1792
rect 13437 1690 13471 1724
rect 13641 1690 13675 1724
rect 13437 1622 13471 1656
rect 13641 1622 13675 1656
rect 13999 2448 14033 2482
rect 13999 2380 14033 2414
rect 13999 2312 14033 2346
rect 13999 2244 14033 2278
rect 13999 2176 14033 2210
rect 13999 2108 14033 2142
rect 13999 2040 14033 2074
rect 13999 1972 14033 2006
rect 13999 1904 14033 1938
rect 13999 1836 14033 1870
rect 13999 1768 14033 1802
rect 13999 1700 14033 1734
rect 13999 1632 14033 1666
rect 13999 1564 14033 1598
rect 14356 2448 14390 2482
rect 14356 2380 14390 2414
rect 14356 2312 14390 2346
rect 14356 2244 14390 2278
rect 14356 2176 14390 2210
rect 14356 2108 14390 2142
rect 14356 2040 14390 2074
rect 14356 1972 14390 2006
rect 14356 1904 14390 1938
rect 14356 1836 14390 1870
rect 14356 1768 14390 1802
rect 14356 1700 14390 1734
rect 14356 1632 14390 1666
rect 14356 1564 14390 1598
<< mvpsubdiff >>
rect 36 5068 15100 5083
rect 36 5049 142 5068
rect 36 5015 51 5049
rect 85 5034 142 5049
rect 176 5034 214 5068
rect 248 5034 286 5068
rect 320 5034 358 5068
rect 392 5034 430 5068
rect 464 5034 502 5068
rect 536 5034 574 5068
rect 608 5034 646 5068
rect 680 5034 718 5068
rect 752 5034 790 5068
rect 824 5034 862 5068
rect 896 5034 934 5068
rect 968 5034 1006 5068
rect 1040 5034 1078 5068
rect 1112 5034 1150 5068
rect 1184 5034 1222 5068
rect 1256 5034 1294 5068
rect 1328 5034 1366 5068
rect 1400 5034 1438 5068
rect 1472 5034 1510 5068
rect 1544 5034 1582 5068
rect 1616 5034 1654 5068
rect 1688 5034 1726 5068
rect 1760 5034 1798 5068
rect 1832 5034 1870 5068
rect 1904 5034 1942 5068
rect 1976 5034 2014 5068
rect 2048 5034 2086 5068
rect 2120 5034 2158 5068
rect 2192 5034 2230 5068
rect 2264 5034 2302 5068
rect 2336 5034 2374 5068
rect 2408 5034 2446 5068
rect 2480 5034 2518 5068
rect 2552 5034 2590 5068
rect 2624 5034 2662 5068
rect 2696 5034 2734 5068
rect 2768 5034 2806 5068
rect 2840 5034 2878 5068
rect 2912 5034 2950 5068
rect 2984 5034 3022 5068
rect 3056 5034 3094 5068
rect 3128 5034 3166 5068
rect 3200 5034 3238 5068
rect 3272 5034 3310 5068
rect 3344 5034 3382 5068
rect 3416 5034 3454 5068
rect 3488 5034 3526 5068
rect 3560 5034 3598 5068
rect 3632 5034 3670 5068
rect 3704 5034 3742 5068
rect 3776 5034 3814 5068
rect 3848 5034 3886 5068
rect 3920 5034 3958 5068
rect 3992 5034 4030 5068
rect 4064 5034 4102 5068
rect 4136 5034 4174 5068
rect 4208 5034 4246 5068
rect 4280 5034 4318 5068
rect 4352 5034 4390 5068
rect 4424 5034 4462 5068
rect 4496 5034 4534 5068
rect 4568 5034 4606 5068
rect 4640 5034 4678 5068
rect 4712 5034 4750 5068
rect 4784 5034 4822 5068
rect 4856 5034 4894 5068
rect 4928 5034 4966 5068
rect 5000 5034 5038 5068
rect 5072 5034 5110 5068
rect 5144 5034 5182 5068
rect 5216 5034 5254 5068
rect 5288 5034 5326 5068
rect 5360 5034 5398 5068
rect 5432 5034 5470 5068
rect 5504 5034 5542 5068
rect 5576 5034 5614 5068
rect 5648 5034 5686 5068
rect 5720 5034 5758 5068
rect 5792 5034 5830 5068
rect 5864 5034 5902 5068
rect 5936 5034 5974 5068
rect 6008 5034 6046 5068
rect 6080 5034 6118 5068
rect 6152 5034 6190 5068
rect 6224 5034 6262 5068
rect 6296 5034 6334 5068
rect 6368 5034 6406 5068
rect 6440 5034 6478 5068
rect 6512 5034 6550 5068
rect 6584 5034 6622 5068
rect 6656 5034 6694 5068
rect 6728 5034 6766 5068
rect 6800 5034 6838 5068
rect 6872 5034 6910 5068
rect 6944 5034 6982 5068
rect 7016 5034 7054 5068
rect 7088 5034 7126 5068
rect 7160 5034 7198 5068
rect 7232 5034 7270 5068
rect 7304 5034 7342 5068
rect 7376 5034 7414 5068
rect 7448 5034 7486 5068
rect 7520 5034 7558 5068
rect 7592 5034 7630 5068
rect 7664 5034 7702 5068
rect 7736 5034 7774 5068
rect 7808 5034 7846 5068
rect 7880 5034 7918 5068
rect 7952 5034 7990 5068
rect 8024 5034 8062 5068
rect 8096 5034 8134 5068
rect 8168 5034 8206 5068
rect 8240 5034 8278 5068
rect 8312 5034 8350 5068
rect 8384 5034 8422 5068
rect 8456 5034 8494 5068
rect 8528 5034 8566 5068
rect 8600 5034 8638 5068
rect 8672 5034 8710 5068
rect 8744 5034 8782 5068
rect 8816 5034 8854 5068
rect 8888 5034 8926 5068
rect 8960 5034 8998 5068
rect 9032 5034 9070 5068
rect 9104 5034 9142 5068
rect 9176 5034 9214 5068
rect 9248 5034 9286 5068
rect 9320 5034 9358 5068
rect 9392 5034 9430 5068
rect 9464 5034 9502 5068
rect 9536 5034 9574 5068
rect 9608 5034 9646 5068
rect 9680 5034 9718 5068
rect 9752 5034 9790 5068
rect 9824 5034 9862 5068
rect 9896 5034 9934 5068
rect 9968 5034 10006 5068
rect 10040 5034 10078 5068
rect 10112 5034 10151 5068
rect 10185 5034 10224 5068
rect 10258 5034 10297 5068
rect 10331 5034 10370 5068
rect 10404 5034 10443 5068
rect 10477 5034 10516 5068
rect 10550 5034 10589 5068
rect 10623 5034 10662 5068
rect 10696 5034 10735 5068
rect 10769 5034 10808 5068
rect 10842 5034 10881 5068
rect 10915 5034 10954 5068
rect 10988 5034 11027 5068
rect 11061 5034 11100 5068
rect 11134 5034 11173 5068
rect 11207 5034 11246 5068
rect 11280 5034 11319 5068
rect 11353 5034 11392 5068
rect 11426 5034 11465 5068
rect 11499 5034 11538 5068
rect 11572 5034 11611 5068
rect 11645 5034 11684 5068
rect 11718 5034 11757 5068
rect 11791 5034 11830 5068
rect 11864 5034 11903 5068
rect 11937 5034 11976 5068
rect 12010 5034 12049 5068
rect 12083 5034 12122 5068
rect 12156 5034 12195 5068
rect 12229 5034 12268 5068
rect 12302 5034 12341 5068
rect 12375 5034 12414 5068
rect 12448 5034 12487 5068
rect 12521 5034 12560 5068
rect 12594 5034 12633 5068
rect 12667 5034 12706 5068
rect 12740 5034 12779 5068
rect 12813 5034 12852 5068
rect 12886 5034 12925 5068
rect 12959 5034 12998 5068
rect 13032 5034 13071 5068
rect 13105 5034 13144 5068
rect 13178 5034 13217 5068
rect 13251 5034 13290 5068
rect 13324 5034 13363 5068
rect 13397 5034 13436 5068
rect 13470 5034 13509 5068
rect 13543 5034 13582 5068
rect 13616 5034 13655 5068
rect 13689 5034 13728 5068
rect 13762 5034 13801 5068
rect 13835 5034 13874 5068
rect 13908 5034 13947 5068
rect 13981 5034 14020 5068
rect 14054 5034 14093 5068
rect 14127 5034 14166 5068
rect 14200 5034 14239 5068
rect 14273 5034 14312 5068
rect 14346 5034 14385 5068
rect 14419 5034 14458 5068
rect 14492 5034 14531 5068
rect 14565 5034 14604 5068
rect 14638 5034 14677 5068
rect 14711 5034 14750 5068
rect 14784 5034 14823 5068
rect 14857 5034 15100 5068
rect 85 5017 15100 5034
rect 85 5015 14915 5017
rect 36 5000 14915 5015
rect 36 4976 119 5000
rect 36 4942 51 4976
rect 85 4966 119 4976
rect 153 4966 191 5000
rect 225 4966 263 5000
rect 297 4966 335 5000
rect 369 4966 407 5000
rect 441 4966 479 5000
rect 513 4966 551 5000
rect 585 4966 623 5000
rect 657 4966 695 5000
rect 729 4966 767 5000
rect 801 4966 839 5000
rect 873 4966 911 5000
rect 945 4966 983 5000
rect 1017 4966 1055 5000
rect 1089 4966 1127 5000
rect 1161 4966 1199 5000
rect 1233 4966 1271 5000
rect 1305 4966 1343 5000
rect 1377 4966 1415 5000
rect 1449 4966 1487 5000
rect 1521 4966 1559 5000
rect 1593 4966 1631 5000
rect 1665 4966 1703 5000
rect 1737 4966 1775 5000
rect 1809 4966 1847 5000
rect 1881 4966 1919 5000
rect 1953 4966 1991 5000
rect 2025 4966 2063 5000
rect 2097 4966 2135 5000
rect 2169 4966 2207 5000
rect 2241 4966 2279 5000
rect 2313 4966 2351 5000
rect 2385 4966 2423 5000
rect 2457 4966 2495 5000
rect 2529 4966 2567 5000
rect 2601 4966 2639 5000
rect 2673 4966 2711 5000
rect 2745 4966 2783 5000
rect 2817 4966 2855 5000
rect 2889 4966 2927 5000
rect 2961 4966 2999 5000
rect 3033 4966 3071 5000
rect 3105 4966 3143 5000
rect 3177 4966 3215 5000
rect 3249 4966 3287 5000
rect 3321 4966 3359 5000
rect 3393 4966 3431 5000
rect 3465 4966 3503 5000
rect 3537 4966 3575 5000
rect 3609 4966 3647 5000
rect 3681 4966 3719 5000
rect 3753 4966 3791 5000
rect 3825 4966 3863 5000
rect 3897 4966 3935 5000
rect 3969 4966 4007 5000
rect 4041 4966 4079 5000
rect 4113 4966 4151 5000
rect 4185 4966 4223 5000
rect 4257 4966 4295 5000
rect 4329 4966 4367 5000
rect 4401 4966 4439 5000
rect 4473 4966 4511 5000
rect 4545 4966 4583 5000
rect 4617 4966 4655 5000
rect 4689 4966 4727 5000
rect 4761 4966 4799 5000
rect 4833 4966 4871 5000
rect 4905 4966 4943 5000
rect 4977 4966 5015 5000
rect 5049 4966 5087 5000
rect 5121 4966 5159 5000
rect 5193 4966 5231 5000
rect 5265 4966 5303 5000
rect 5337 4966 5375 5000
rect 5409 4966 5447 5000
rect 5481 4966 5519 5000
rect 5553 4966 5591 5000
rect 5625 4966 5663 5000
rect 5697 4966 5735 5000
rect 5769 4966 5807 5000
rect 5841 4966 5879 5000
rect 5913 4966 5951 5000
rect 5985 4966 6023 5000
rect 6057 4966 6095 5000
rect 6129 4966 6167 5000
rect 6201 4966 6239 5000
rect 6273 4966 6311 5000
rect 6345 4966 6383 5000
rect 6417 4966 6455 5000
rect 6489 4966 6527 5000
rect 6561 4966 6599 5000
rect 6633 4966 6671 5000
rect 6705 4966 6743 5000
rect 6777 4966 6815 5000
rect 6849 4966 6887 5000
rect 6921 4966 6959 5000
rect 6993 4966 7031 5000
rect 7065 4966 7103 5000
rect 7137 4966 7175 5000
rect 7209 4966 7247 5000
rect 7281 4966 7319 5000
rect 7353 4966 7391 5000
rect 7425 4966 7463 5000
rect 7497 4966 7535 5000
rect 7569 4966 7607 5000
rect 7641 4966 7679 5000
rect 7713 4966 7751 5000
rect 7785 4966 7823 5000
rect 7857 4966 7895 5000
rect 7929 4966 7967 5000
rect 8001 4966 8039 5000
rect 8073 4966 8111 5000
rect 8145 4966 8183 5000
rect 8217 4966 8255 5000
rect 8289 4966 8327 5000
rect 8361 4966 8399 5000
rect 8433 4966 8471 5000
rect 8505 4966 8543 5000
rect 8577 4966 8615 5000
rect 8649 4966 8687 5000
rect 8721 4966 8759 5000
rect 8793 4966 8831 5000
rect 8865 4966 8903 5000
rect 8937 4966 8975 5000
rect 9009 4966 9047 5000
rect 9081 4966 9119 5000
rect 9153 4966 9191 5000
rect 9225 4966 9263 5000
rect 9297 4966 9335 5000
rect 9369 4966 9407 5000
rect 9441 4966 9479 5000
rect 9513 4966 9551 5000
rect 9585 4966 9623 5000
rect 9657 4966 9695 5000
rect 9729 4966 9767 5000
rect 9801 4966 9839 5000
rect 9873 4966 9911 5000
rect 9945 4966 9983 5000
rect 10017 4966 10055 5000
rect 10089 4966 10127 5000
rect 10161 4966 10199 5000
rect 10233 4966 10271 5000
rect 10305 4966 10343 5000
rect 10377 4966 10415 5000
rect 10449 4966 10487 5000
rect 10521 4966 10559 5000
rect 10593 4966 10631 5000
rect 10665 4966 10703 5000
rect 10737 4966 10775 5000
rect 10809 4966 10847 5000
rect 10881 4966 10919 5000
rect 10953 4966 10991 5000
rect 11025 4966 11063 5000
rect 11097 4966 11135 5000
rect 11169 4966 11207 5000
rect 11241 4966 11279 5000
rect 11313 4966 11351 5000
rect 11385 4966 11423 5000
rect 11457 4966 11495 5000
rect 11529 4966 11567 5000
rect 11601 4966 11639 5000
rect 11673 4966 11711 5000
rect 11745 4966 11783 5000
rect 11817 4966 11855 5000
rect 11889 4966 11927 5000
rect 11961 4966 11999 5000
rect 12033 4966 12071 5000
rect 12105 4966 12143 5000
rect 12177 4966 12215 5000
rect 12249 4966 12287 5000
rect 12321 4966 12359 5000
rect 12393 4966 12431 5000
rect 12465 4966 12503 5000
rect 12537 4966 12575 5000
rect 12609 4966 12647 5000
rect 12681 4966 12719 5000
rect 12753 4966 12791 5000
rect 12825 4966 12863 5000
rect 12897 4966 12935 5000
rect 12969 4966 13007 5000
rect 13041 4966 13079 5000
rect 13113 4966 13151 5000
rect 13185 4966 13223 5000
rect 13257 4966 13295 5000
rect 13329 4966 13367 5000
rect 13401 4966 13439 5000
rect 13473 4966 13511 5000
rect 13545 4966 13583 5000
rect 13617 4966 13655 5000
rect 13689 4966 13728 5000
rect 13762 4966 13801 5000
rect 13835 4966 13874 5000
rect 13908 4966 13947 5000
rect 13981 4966 14020 5000
rect 14054 4966 14093 5000
rect 14127 4966 14166 5000
rect 14200 4966 14239 5000
rect 14273 4966 14312 5000
rect 14346 4966 14385 5000
rect 14419 4966 14458 5000
rect 14492 4966 14531 5000
rect 14565 4966 14604 5000
rect 14638 4966 14677 5000
rect 14711 4966 14750 5000
rect 14784 4966 14823 5000
rect 14857 4983 14915 5000
rect 14949 4983 14983 5017
rect 15017 4983 15051 5017
rect 15085 4983 15100 5017
rect 14857 4966 15100 4983
rect 85 4945 15100 4966
rect 85 4942 14915 4945
rect 36 4932 14915 4942
rect 36 4926 187 4932
rect 36 4903 119 4926
rect 36 4869 51 4903
rect 85 4892 119 4903
rect 153 4898 187 4926
rect 221 4898 259 4932
rect 293 4898 331 4932
rect 365 4898 403 4932
rect 437 4898 475 4932
rect 509 4898 547 4932
rect 581 4898 619 4932
rect 653 4898 691 4932
rect 725 4898 763 4932
rect 797 4898 835 4932
rect 869 4898 907 4932
rect 941 4898 979 4932
rect 1013 4898 1051 4932
rect 1085 4898 1123 4932
rect 1157 4898 1195 4932
rect 1229 4898 1267 4932
rect 1301 4898 1339 4932
rect 1373 4898 1411 4932
rect 1445 4898 1483 4932
rect 1517 4898 1555 4932
rect 1589 4898 1627 4932
rect 1661 4898 1699 4932
rect 1733 4898 1771 4932
rect 1805 4898 1843 4932
rect 1877 4898 1915 4932
rect 1949 4898 1987 4932
rect 2021 4898 2059 4932
rect 2093 4898 2131 4932
rect 2165 4898 2203 4932
rect 2237 4898 2275 4932
rect 2309 4898 2347 4932
rect 2381 4898 2419 4932
rect 2453 4898 2491 4932
rect 2525 4898 2563 4932
rect 2597 4898 2635 4932
rect 2669 4898 2707 4932
rect 2741 4898 2779 4932
rect 2813 4898 2851 4932
rect 2885 4898 2923 4932
rect 2957 4898 2995 4932
rect 3029 4898 3067 4932
rect 3101 4898 3139 4932
rect 3173 4898 3211 4932
rect 3245 4898 3283 4932
rect 3317 4898 3355 4932
rect 3389 4898 3427 4932
rect 3461 4898 3499 4932
rect 3533 4898 3571 4932
rect 3605 4898 3643 4932
rect 3677 4898 3715 4932
rect 3749 4898 3787 4932
rect 3821 4898 3859 4932
rect 3893 4898 3931 4932
rect 3965 4898 4003 4932
rect 4037 4898 4075 4932
rect 4109 4898 4147 4932
rect 4181 4898 4219 4932
rect 4253 4898 4291 4932
rect 4325 4898 4363 4932
rect 4397 4898 4435 4932
rect 4469 4898 4507 4932
rect 4541 4898 4579 4932
rect 4613 4898 4651 4932
rect 4685 4898 4723 4932
rect 4757 4898 4795 4932
rect 4829 4898 4867 4932
rect 4901 4898 4939 4932
rect 4973 4898 5011 4932
rect 5045 4898 5083 4932
rect 5117 4898 5155 4932
rect 5189 4898 5227 4932
rect 5261 4898 5299 4932
rect 5333 4898 5371 4932
rect 5405 4898 5443 4932
rect 5477 4898 5515 4932
rect 5549 4898 5587 4932
rect 5621 4898 5659 4932
rect 5693 4898 5731 4932
rect 5765 4898 5803 4932
rect 5837 4898 5875 4932
rect 5909 4898 5947 4932
rect 5981 4898 6019 4932
rect 6053 4898 6091 4932
rect 6125 4898 6163 4932
rect 6197 4898 6235 4932
rect 6269 4898 6307 4932
rect 6341 4898 6379 4932
rect 6413 4898 6451 4932
rect 6485 4898 6523 4932
rect 6557 4898 6595 4932
rect 6629 4898 6667 4932
rect 6701 4898 6739 4932
rect 6773 4898 6811 4932
rect 6845 4898 6883 4932
rect 6917 4898 6955 4932
rect 6989 4898 7027 4932
rect 7061 4898 7099 4932
rect 7133 4898 7171 4932
rect 7205 4898 7243 4932
rect 7277 4898 7315 4932
rect 7349 4898 7387 4932
rect 7421 4898 7459 4932
rect 7493 4898 7531 4932
rect 7565 4898 7603 4932
rect 7637 4898 7675 4932
rect 7709 4898 7747 4932
rect 7781 4898 7819 4932
rect 7853 4898 7891 4932
rect 7925 4898 7963 4932
rect 7997 4898 8035 4932
rect 8069 4898 8107 4932
rect 8141 4898 8179 4932
rect 8213 4898 8251 4932
rect 8285 4898 8323 4932
rect 8357 4898 8395 4932
rect 8429 4898 8467 4932
rect 8501 4898 8539 4932
rect 8573 4898 8611 4932
rect 8645 4898 8683 4932
rect 8717 4898 8755 4932
rect 8789 4898 8827 4932
rect 8861 4898 8899 4932
rect 8933 4898 8971 4932
rect 9005 4898 9043 4932
rect 9077 4898 9115 4932
rect 9149 4898 9187 4932
rect 9221 4898 9259 4932
rect 9293 4898 9331 4932
rect 9365 4898 9403 4932
rect 9437 4898 9475 4932
rect 9509 4898 9547 4932
rect 9581 4898 9619 4932
rect 9653 4898 9691 4932
rect 9725 4898 9763 4932
rect 9797 4898 9835 4932
rect 9869 4898 9907 4932
rect 9941 4898 9979 4932
rect 10013 4898 10051 4932
rect 10085 4898 10123 4932
rect 10157 4898 10195 4932
rect 10229 4898 10267 4932
rect 10301 4898 10339 4932
rect 10373 4898 10411 4932
rect 10445 4898 10483 4932
rect 10517 4898 10555 4932
rect 10589 4898 10627 4932
rect 10661 4898 10699 4932
rect 10733 4898 10771 4932
rect 10805 4898 10843 4932
rect 10877 4898 10915 4932
rect 10949 4898 10987 4932
rect 11021 4898 11059 4932
rect 11093 4898 11131 4932
rect 11165 4898 11203 4932
rect 11237 4898 11275 4932
rect 11309 4898 11347 4932
rect 11381 4898 11419 4932
rect 11453 4898 11491 4932
rect 11525 4898 11563 4932
rect 11597 4898 11635 4932
rect 11669 4898 11707 4932
rect 11741 4898 11779 4932
rect 11813 4898 11851 4932
rect 11885 4898 11923 4932
rect 11957 4898 11995 4932
rect 12029 4898 12067 4932
rect 12101 4898 12139 4932
rect 12173 4898 12211 4932
rect 12245 4898 12283 4932
rect 12317 4898 12355 4932
rect 12389 4898 12427 4932
rect 12461 4898 12499 4932
rect 12533 4898 12571 4932
rect 12605 4898 12643 4932
rect 12677 4898 12715 4932
rect 12749 4898 12787 4932
rect 12821 4898 12859 4932
rect 12893 4898 12931 4932
rect 12965 4898 13003 4932
rect 13037 4898 13075 4932
rect 13109 4898 13147 4932
rect 13181 4898 13219 4932
rect 13253 4898 13291 4932
rect 13325 4898 13363 4932
rect 13397 4898 13436 4932
rect 13470 4898 13509 4932
rect 13543 4898 13582 4932
rect 13616 4898 13655 4932
rect 13689 4898 13728 4932
rect 13762 4898 13801 4932
rect 13835 4898 13874 4932
rect 13908 4898 13947 4932
rect 13981 4898 14020 4932
rect 14054 4898 14093 4932
rect 14127 4898 14166 4932
rect 14200 4898 14239 4932
rect 14273 4898 14312 4932
rect 14346 4898 14385 4932
rect 14419 4898 14458 4932
rect 14492 4898 14531 4932
rect 14565 4898 14604 4932
rect 14638 4898 14677 4932
rect 14711 4898 14750 4932
rect 14784 4898 14823 4932
rect 14857 4911 14915 4932
rect 14949 4911 14983 4945
rect 15017 4911 15051 4945
rect 15085 4911 15100 4945
rect 14857 4898 15100 4911
rect 153 4892 15100 4898
rect 85 4883 15100 4892
rect 85 4869 329 4883
rect 36 4859 329 4869
rect 36 4857 262 4859
rect 36 4852 187 4857
rect 36 4830 119 4852
rect 36 4796 51 4830
rect 85 4818 119 4830
rect 153 4823 187 4852
rect 221 4825 262 4857
rect 296 4825 329 4859
rect 221 4823 329 4825
rect 153 4818 329 4823
rect 85 4796 329 4818
rect 36 4791 329 4796
rect 36 4782 262 4791
rect 36 4778 187 4782
rect 36 4757 119 4778
rect 36 4723 51 4757
rect 85 4744 119 4757
rect 153 4748 187 4778
rect 221 4757 262 4782
rect 296 4757 329 4791
rect 221 4748 329 4757
rect 153 4744 329 4748
rect 85 4723 329 4744
rect 36 4707 262 4723
rect 36 4704 187 4707
rect 36 4684 119 4704
rect 36 4650 51 4684
rect 85 4670 119 4684
rect 153 4673 187 4704
rect 221 4689 262 4707
rect 296 4689 329 4723
rect 221 4673 329 4689
rect 153 4670 329 4673
rect 85 4655 329 4670
rect 85 4650 262 4655
rect 36 4632 262 4650
rect 36 4630 187 4632
rect 36 4611 119 4630
rect 36 4577 51 4611
rect 85 4596 119 4611
rect 153 4598 187 4630
rect 221 4621 262 4632
rect 296 4621 329 4655
rect 14807 4873 15100 4883
rect 14807 4859 14915 4873
rect 14807 4825 14840 4859
rect 14874 4839 14915 4859
rect 14949 4839 14983 4873
rect 15017 4839 15051 4873
rect 15085 4839 15100 4873
rect 14874 4825 15100 4839
rect 14807 4801 15100 4825
rect 14807 4791 14915 4801
rect 14807 4757 14840 4791
rect 14874 4767 14915 4791
rect 14949 4767 14983 4801
rect 15017 4767 15051 4801
rect 15085 4767 15100 4801
rect 14874 4757 15100 4767
rect 14807 4729 15100 4757
rect 14807 4723 14915 4729
rect 14807 4689 14840 4723
rect 14874 4695 14915 4723
rect 14949 4695 14983 4729
rect 15017 4695 15051 4729
rect 15085 4695 15100 4729
rect 14874 4689 15100 4695
rect 14807 4657 15100 4689
rect 14807 4655 14915 4657
rect 221 4598 329 4621
rect 153 4596 329 4598
rect 85 4587 329 4596
rect 85 4577 262 4587
rect 36 4557 262 4577
rect 36 4556 187 4557
rect 36 4538 119 4556
rect 36 4504 51 4538
rect 85 4522 119 4538
rect 153 4523 187 4556
rect 221 4553 262 4557
rect 296 4553 329 4587
rect 221 4523 329 4553
rect 153 4522 329 4523
rect 85 4519 329 4522
rect 85 4504 262 4519
rect 36 4485 262 4504
rect 296 4485 329 4519
rect 36 4483 329 4485
rect 36 4482 187 4483
rect 36 4465 119 4482
rect 36 4431 51 4465
rect 85 4448 119 4465
rect 153 4449 187 4482
rect 221 4451 329 4483
rect 221 4449 262 4451
rect 153 4448 262 4449
rect 85 4431 262 4448
rect 36 4417 262 4431
rect 296 4417 329 4451
rect 36 4409 329 4417
rect 36 4408 187 4409
rect 36 4393 119 4408
rect 36 4359 51 4393
rect 85 4374 119 4393
rect 153 4375 187 4408
rect 221 4383 329 4409
rect 221 4375 262 4383
rect 153 4374 262 4375
rect 85 4359 262 4374
rect 36 4349 262 4359
rect 296 4349 329 4383
rect 36 4335 329 4349
rect 36 4334 187 4335
rect 36 4321 119 4334
rect 36 4287 51 4321
rect 85 4300 119 4321
rect 153 4301 187 4334
rect 221 4315 329 4335
rect 221 4301 262 4315
rect 153 4300 262 4301
rect 85 4287 262 4300
rect 36 4281 262 4287
rect 296 4281 329 4315
rect 36 4261 329 4281
rect 36 4260 187 4261
rect 36 4249 119 4260
rect 36 4215 51 4249
rect 85 4226 119 4249
rect 153 4227 187 4260
rect 221 4247 329 4261
rect 221 4227 262 4247
rect 153 4226 262 4227
rect 85 4215 262 4226
rect 36 4213 262 4215
rect 296 4213 329 4247
rect 36 4187 329 4213
rect 36 4186 187 4187
rect 36 4177 119 4186
rect 36 4143 51 4177
rect 85 4152 119 4177
rect 153 4153 187 4186
rect 221 4179 329 4187
rect 221 4153 262 4179
rect 153 4152 262 4153
rect 85 4145 262 4152
rect 296 4145 329 4179
rect 85 4143 329 4145
rect 36 4113 329 4143
rect 36 4112 187 4113
rect 36 4105 119 4112
rect 36 4071 51 4105
rect 85 4078 119 4105
rect 153 4079 187 4112
rect 221 4111 329 4113
rect 221 4079 262 4111
rect 153 4078 262 4079
rect 85 4077 262 4078
rect 296 4077 329 4111
rect 85 4071 329 4077
rect 36 4043 329 4071
rect 36 4039 262 4043
rect 36 4038 187 4039
rect 36 4033 119 4038
rect 36 3999 51 4033
rect 85 4004 119 4033
rect 153 4005 187 4038
rect 221 4009 262 4039
rect 296 4009 329 4043
rect 221 4005 329 4009
rect 153 4004 329 4005
rect 85 3999 329 4004
rect 36 3975 329 3999
rect 36 3965 262 3975
rect 36 3964 187 3965
rect 36 3961 119 3964
rect 36 3927 51 3961
rect 85 3930 119 3961
rect 153 3931 187 3964
rect 221 3941 262 3965
rect 296 3941 329 3975
rect 221 3931 329 3941
rect 153 3930 329 3931
rect 85 3927 329 3930
rect 36 3907 329 3927
rect 36 3891 262 3907
rect 36 3890 187 3891
rect 36 3889 119 3890
rect 36 3855 51 3889
rect 85 3856 119 3889
rect 153 3857 187 3890
rect 221 3873 262 3891
rect 296 3873 329 3907
rect 221 3857 329 3873
rect 153 3856 329 3857
rect 85 3855 329 3856
rect 36 3839 329 3855
rect 36 3817 262 3839
rect 36 3783 51 3817
rect 85 3783 119 3817
rect 153 3783 187 3817
rect 221 3805 262 3817
rect 296 3805 329 3839
rect 221 3783 329 3805
rect 36 3771 329 3783
rect 36 3737 262 3771
rect 296 3737 329 3771
rect 36 3707 329 3737
rect 36 3673 51 3707
rect 85 3673 119 3707
rect 153 3673 187 3707
rect 221 3703 329 3707
rect 221 3673 262 3703
rect 36 3669 262 3673
rect 296 3669 329 3703
rect 36 3635 329 3669
rect 36 3634 262 3635
rect 36 3600 51 3634
rect 85 3600 119 3634
rect 153 3600 187 3634
rect 221 3601 262 3634
rect 296 3601 329 3635
rect 221 3600 329 3601
rect 36 3567 329 3600
rect 36 3562 262 3567
rect 36 3528 51 3562
rect 85 3528 119 3562
rect 153 3528 187 3562
rect 221 3533 262 3562
rect 296 3533 329 3567
rect 221 3528 329 3533
rect 36 3499 329 3528
rect 36 3490 262 3499
rect 36 3456 51 3490
rect 85 3456 119 3490
rect 153 3456 187 3490
rect 221 3465 262 3490
rect 296 3465 329 3499
rect 221 3456 329 3465
rect 36 3431 329 3456
rect 36 3418 262 3431
rect 36 3384 51 3418
rect 85 3384 119 3418
rect 153 3384 187 3418
rect 221 3397 262 3418
rect 296 3397 329 3431
rect 221 3384 329 3397
rect 36 3363 329 3384
rect 36 3346 262 3363
rect 36 3312 51 3346
rect 85 3312 119 3346
rect 153 3312 187 3346
rect 221 3329 262 3346
rect 296 3329 329 3363
rect 221 3312 329 3329
rect 36 3295 329 3312
rect 36 3274 262 3295
rect 36 3240 51 3274
rect 85 3240 119 3274
rect 153 3240 187 3274
rect 221 3261 262 3274
rect 296 3261 329 3295
rect 221 3240 329 3261
rect 36 3227 329 3240
rect 36 3202 262 3227
rect 36 3168 51 3202
rect 85 3168 119 3202
rect 153 3168 187 3202
rect 221 3193 262 3202
rect 296 3193 329 3227
rect 221 3168 329 3193
rect 36 3159 329 3168
rect 36 3130 262 3159
rect 36 3096 51 3130
rect 85 3096 119 3130
rect 153 3096 187 3130
rect 221 3125 262 3130
rect 296 3125 329 3159
rect 221 3096 329 3125
rect 36 3091 329 3096
rect 36 3058 262 3091
rect 36 3024 51 3058
rect 85 3024 119 3058
rect 153 3024 187 3058
rect 221 3057 262 3058
rect 296 3057 329 3091
rect 221 3024 329 3057
rect 36 3023 329 3024
rect 36 2989 262 3023
rect 296 2989 329 3023
rect 36 2986 329 2989
rect 36 2952 51 2986
rect 85 2952 119 2986
rect 153 2952 187 2986
rect 221 2955 329 2986
rect 221 2952 262 2955
rect 36 2921 262 2952
rect 296 2921 329 2955
rect 36 2914 329 2921
rect 36 2880 51 2914
rect 85 2880 119 2914
rect 153 2880 187 2914
rect 221 2887 329 2914
rect 221 2880 262 2887
rect 36 2853 262 2880
rect 296 2853 329 2887
rect 36 2842 329 2853
rect 36 2808 51 2842
rect 85 2808 119 2842
rect 153 2808 187 2842
rect 221 2819 329 2842
rect 221 2808 262 2819
rect 36 2785 262 2808
rect 296 2785 329 2819
rect 36 2770 329 2785
rect 36 2736 51 2770
rect 85 2736 119 2770
rect 153 2736 187 2770
rect 221 2751 329 2770
rect 221 2736 262 2751
rect 36 2717 262 2736
rect 296 2717 329 2751
rect 36 2698 329 2717
rect 36 2664 51 2698
rect 85 2664 119 2698
rect 153 2664 187 2698
rect 221 2683 329 2698
rect 221 2664 262 2683
rect 36 2649 262 2664
rect 296 2649 329 2683
rect 36 2626 329 2649
rect 36 2592 51 2626
rect 85 2592 119 2626
rect 153 2592 187 2626
rect 221 2615 329 2626
rect 221 2592 262 2615
rect 36 2581 262 2592
rect 296 2581 329 2615
rect 36 2554 329 2581
rect 36 2520 51 2554
rect 85 2520 119 2554
rect 153 2520 187 2554
rect 221 2547 329 2554
rect 221 2520 262 2547
rect 36 2513 262 2520
rect 296 2513 329 2547
rect 36 2482 329 2513
rect 36 2448 51 2482
rect 85 2448 119 2482
rect 153 2448 187 2482
rect 221 2479 329 2482
rect 221 2448 262 2479
rect 36 2445 262 2448
rect 296 2445 329 2479
rect 36 2411 329 2445
rect 36 2410 262 2411
rect 36 2376 51 2410
rect 85 2376 119 2410
rect 153 2376 187 2410
rect 221 2377 262 2410
rect 296 2377 329 2411
rect 221 2376 329 2377
rect 36 2343 329 2376
rect 36 2338 262 2343
rect 36 2304 51 2338
rect 85 2304 119 2338
rect 153 2304 187 2338
rect 221 2309 262 2338
rect 296 2309 329 2343
rect 221 2304 329 2309
rect 36 2275 329 2304
rect 36 2266 262 2275
rect 36 2232 51 2266
rect 85 2232 119 2266
rect 153 2232 187 2266
rect 221 2241 262 2266
rect 296 2241 329 2275
rect 221 2232 329 2241
rect 36 2207 329 2232
rect 36 2194 262 2207
rect 36 2160 51 2194
rect 85 2160 119 2194
rect 153 2160 187 2194
rect 221 2173 262 2194
rect 296 2173 329 2207
rect 221 2160 329 2173
rect 36 2139 329 2160
rect 36 2122 262 2139
rect 36 2088 51 2122
rect 85 2088 119 2122
rect 153 2088 187 2122
rect 221 2105 262 2122
rect 296 2105 329 2139
rect 221 2088 329 2105
rect 36 2071 329 2088
rect 36 2050 262 2071
rect 36 2016 51 2050
rect 85 2016 119 2050
rect 153 2016 187 2050
rect 221 2037 262 2050
rect 296 2037 329 2071
rect 221 2016 329 2037
rect 36 2003 329 2016
rect 36 1978 262 2003
rect 36 1944 51 1978
rect 85 1944 119 1978
rect 153 1944 187 1978
rect 221 1969 262 1978
rect 296 1969 329 2003
rect 221 1944 329 1969
rect 36 1935 329 1944
rect 36 1906 262 1935
rect 36 1872 51 1906
rect 85 1872 119 1906
rect 153 1872 187 1906
rect 221 1901 262 1906
rect 296 1901 329 1935
rect 221 1872 329 1901
rect 36 1867 329 1872
rect 36 1834 262 1867
rect 36 1800 51 1834
rect 85 1800 119 1834
rect 153 1800 187 1834
rect 221 1833 262 1834
rect 296 1833 329 1867
rect 221 1800 329 1833
rect 36 1799 329 1800
rect 36 1765 262 1799
rect 296 1765 329 1799
rect 36 1762 329 1765
rect 36 1728 51 1762
rect 85 1728 119 1762
rect 153 1728 187 1762
rect 221 1731 329 1762
rect 221 1728 262 1731
rect 36 1697 262 1728
rect 296 1697 329 1731
rect 36 1690 329 1697
rect 36 1656 51 1690
rect 85 1656 119 1690
rect 153 1656 187 1690
rect 221 1663 329 1690
rect 221 1656 262 1663
rect 36 1629 262 1656
rect 296 1629 329 1663
rect 36 1618 329 1629
rect 36 1584 51 1618
rect 85 1584 119 1618
rect 153 1584 187 1618
rect 221 1595 329 1618
rect 221 1584 262 1595
rect 36 1561 262 1584
rect 296 1561 329 1595
rect 36 1546 329 1561
rect 36 1512 51 1546
rect 85 1512 119 1546
rect 153 1512 187 1546
rect 221 1527 329 1546
rect 221 1512 262 1527
rect 36 1493 262 1512
rect 296 1493 329 1527
rect 36 1474 329 1493
rect 36 1440 51 1474
rect 85 1440 119 1474
rect 153 1440 187 1474
rect 221 1459 329 1474
rect 221 1440 262 1459
rect 36 1425 262 1440
rect 296 1425 329 1459
rect 36 1402 329 1425
rect 36 1368 51 1402
rect 85 1368 119 1402
rect 153 1368 187 1402
rect 221 1391 329 1402
rect 221 1368 262 1391
rect 36 1357 262 1368
rect 296 1357 329 1391
rect 36 1330 329 1357
rect 36 1296 51 1330
rect 85 1296 119 1330
rect 153 1296 187 1330
rect 221 1323 329 1330
rect 221 1296 262 1323
rect 36 1289 262 1296
rect 296 1289 329 1323
rect 36 1258 329 1289
rect 36 1224 51 1258
rect 85 1224 119 1258
rect 153 1224 187 1258
rect 221 1255 329 1258
rect 221 1224 262 1255
rect 36 1221 262 1224
rect 296 1221 329 1255
rect 36 1187 329 1221
rect 36 1186 262 1187
rect 36 1152 51 1186
rect 85 1152 119 1186
rect 153 1152 187 1186
rect 221 1153 262 1186
rect 296 1153 329 1187
rect 221 1152 329 1153
rect 36 1119 329 1152
rect 36 1114 262 1119
rect 36 1080 51 1114
rect 85 1080 119 1114
rect 153 1080 187 1114
rect 221 1085 262 1114
rect 296 1085 329 1119
rect 221 1080 329 1085
rect 36 1051 329 1080
rect 36 1042 262 1051
rect 36 1008 51 1042
rect 85 1008 119 1042
rect 153 1008 187 1042
rect 221 1017 262 1042
rect 296 1017 329 1051
rect 221 1008 329 1017
rect 36 983 329 1008
rect 36 970 262 983
rect 36 936 51 970
rect 85 936 119 970
rect 153 936 187 970
rect 221 949 262 970
rect 296 949 329 983
rect 221 936 329 949
rect 36 915 329 936
rect 36 898 262 915
rect 36 864 51 898
rect 85 864 119 898
rect 153 864 187 898
rect 221 881 262 898
rect 296 881 329 915
rect 221 864 329 881
rect 36 847 329 864
rect 36 826 262 847
rect 36 792 51 826
rect 85 792 119 826
rect 153 792 187 826
rect 221 813 262 826
rect 296 813 329 847
rect 221 792 329 813
rect 36 779 329 792
rect 36 754 262 779
rect 36 720 51 754
rect 85 720 119 754
rect 153 720 187 754
rect 221 745 262 754
rect 296 745 329 779
rect 221 720 329 745
rect 36 711 329 720
rect 36 682 262 711
rect 36 648 51 682
rect 85 648 119 682
rect 153 648 187 682
rect 221 677 262 682
rect 296 677 329 711
rect 221 648 329 677
rect 14807 4621 14840 4655
rect 14874 4623 14915 4655
rect 14949 4623 14983 4657
rect 15017 4623 15051 4657
rect 15085 4623 15100 4657
rect 14874 4621 15100 4623
rect 14807 4587 15100 4621
rect 14807 4553 14840 4587
rect 14874 4585 15100 4587
rect 14874 4553 14915 4585
rect 14807 4551 14915 4553
rect 14949 4551 14983 4585
rect 15017 4551 15051 4585
rect 15085 4551 15100 4585
rect 14807 4519 15100 4551
rect 14807 4485 14840 4519
rect 14874 4513 15100 4519
rect 14874 4485 14915 4513
rect 14807 4479 14915 4485
rect 14949 4479 14983 4513
rect 15017 4479 15051 4513
rect 15085 4479 15100 4513
rect 14807 4451 15100 4479
rect 14807 4417 14840 4451
rect 14874 4441 15100 4451
rect 14874 4417 14915 4441
rect 14807 4407 14915 4417
rect 14949 4407 14983 4441
rect 15017 4407 15051 4441
rect 15085 4407 15100 4441
rect 14807 4383 15100 4407
rect 14807 4349 14840 4383
rect 14874 4369 15100 4383
rect 14874 4368 14983 4369
rect 14874 4349 14915 4368
rect 14807 4334 14915 4349
rect 14949 4335 14983 4368
rect 15017 4335 15051 4369
rect 15085 4335 15100 4369
rect 14949 4334 15100 4335
rect 14807 4315 15100 4334
rect 14807 4281 14840 4315
rect 14874 4297 15100 4315
rect 14874 4295 14983 4297
rect 14874 4281 14915 4295
rect 14807 4261 14915 4281
rect 14949 4263 14983 4295
rect 15017 4263 15051 4297
rect 15085 4263 15100 4297
rect 14949 4261 15100 4263
rect 14807 4247 15100 4261
rect 14807 4213 14840 4247
rect 14874 4225 15100 4247
rect 14874 4222 14983 4225
rect 14874 4213 14915 4222
rect 14807 4188 14915 4213
rect 14949 4191 14983 4222
rect 15017 4191 15051 4225
rect 15085 4191 15100 4225
rect 14949 4188 15100 4191
rect 14807 4179 15100 4188
rect 14807 4145 14840 4179
rect 14874 4153 15100 4179
rect 14874 4149 14983 4153
rect 14874 4145 14915 4149
rect 14807 4115 14915 4145
rect 14949 4119 14983 4149
rect 15017 4119 15051 4153
rect 15085 4119 15100 4153
rect 14949 4115 15100 4119
rect 14807 4111 15100 4115
rect 14807 4077 14840 4111
rect 14874 4081 15100 4111
rect 14874 4077 14983 4081
rect 14807 4076 14983 4077
rect 14807 4043 14915 4076
rect 14807 4009 14840 4043
rect 14874 4042 14915 4043
rect 14949 4047 14983 4076
rect 15017 4047 15051 4081
rect 15085 4047 15100 4081
rect 14949 4042 15100 4047
rect 14874 4009 15100 4042
rect 14807 4008 15051 4009
rect 14807 4003 14983 4008
rect 14807 3975 14915 4003
rect 14807 3941 14840 3975
rect 14874 3969 14915 3975
rect 14949 3974 14983 4003
rect 15017 3975 15051 4008
rect 15085 3975 15100 4009
rect 15017 3974 15100 3975
rect 14949 3969 15100 3974
rect 14874 3941 15100 3969
rect 14807 3937 15100 3941
rect 14807 3935 15051 3937
rect 14807 3930 14983 3935
rect 14807 3907 14915 3930
rect 14807 3873 14840 3907
rect 14874 3896 14915 3907
rect 14949 3901 14983 3930
rect 15017 3903 15051 3935
rect 15085 3903 15100 3937
rect 15017 3901 15100 3903
rect 14949 3896 15100 3901
rect 14874 3873 15100 3896
rect 14807 3865 15100 3873
rect 14807 3862 15051 3865
rect 14807 3857 14983 3862
rect 14807 3839 14915 3857
rect 14807 3805 14840 3839
rect 14874 3823 14915 3839
rect 14949 3828 14983 3857
rect 15017 3831 15051 3862
rect 15085 3831 15100 3865
rect 15017 3828 15100 3831
rect 14949 3823 15100 3828
rect 14874 3805 15100 3823
rect 14807 3793 15100 3805
rect 14807 3789 15051 3793
rect 14807 3784 14983 3789
rect 14807 3771 14915 3784
rect 14807 3737 14840 3771
rect 14874 3750 14915 3771
rect 14949 3755 14983 3784
rect 15017 3759 15051 3789
rect 15085 3759 15100 3793
rect 15017 3755 15100 3759
rect 14949 3750 15100 3755
rect 14874 3737 15100 3750
rect 14807 3721 15100 3737
rect 14807 3716 15051 3721
rect 14807 3711 14983 3716
rect 14807 3703 14915 3711
rect 14807 3669 14840 3703
rect 14874 3677 14915 3703
rect 14949 3682 14983 3711
rect 15017 3687 15051 3716
rect 15085 3687 15100 3721
rect 15017 3682 15100 3687
rect 14949 3677 15100 3682
rect 14874 3669 15100 3677
rect 14807 3649 15100 3669
rect 14807 3643 15051 3649
rect 14807 3638 14983 3643
rect 14807 3635 14915 3638
rect 14807 3601 14840 3635
rect 14874 3604 14915 3635
rect 14949 3609 14983 3638
rect 15017 3615 15051 3643
rect 15085 3615 15100 3649
rect 15017 3609 15100 3615
rect 14949 3604 15100 3609
rect 14874 3601 15100 3604
rect 14807 3577 15100 3601
rect 14807 3570 15051 3577
rect 14807 3567 14983 3570
rect 14807 3533 14840 3567
rect 14874 3565 14983 3567
rect 14874 3533 14915 3565
rect 14807 3531 14915 3533
rect 14949 3536 14983 3565
rect 15017 3543 15051 3570
rect 15085 3543 15100 3577
rect 15017 3536 15100 3543
rect 14949 3531 15100 3536
rect 14807 3505 15100 3531
rect 14807 3499 15051 3505
rect 14807 3465 14840 3499
rect 14874 3497 15051 3499
rect 14874 3492 14983 3497
rect 14874 3465 14915 3492
rect 14807 3458 14915 3465
rect 14949 3463 14983 3492
rect 15017 3471 15051 3497
rect 15085 3471 15100 3505
rect 15017 3463 15100 3471
rect 14949 3458 15100 3463
rect 14807 3433 15100 3458
rect 14807 3431 15051 3433
rect 14807 3397 14840 3431
rect 14874 3424 15051 3431
rect 14874 3419 14983 3424
rect 14874 3397 14915 3419
rect 14807 3385 14915 3397
rect 14949 3390 14983 3419
rect 15017 3399 15051 3424
rect 15085 3399 15100 3433
rect 15017 3390 15100 3399
rect 14949 3385 15100 3390
rect 14807 3363 15100 3385
rect 14807 3329 14840 3363
rect 14874 3361 15100 3363
rect 14874 3351 15051 3361
rect 14874 3346 14983 3351
rect 14874 3329 14915 3346
rect 14807 3312 14915 3329
rect 14949 3317 14983 3346
rect 15017 3327 15051 3351
rect 15085 3327 15100 3361
rect 15017 3317 15100 3327
rect 14949 3312 15100 3317
rect 14807 3295 15100 3312
rect 14807 3261 14840 3295
rect 14874 3289 15100 3295
rect 14874 3278 15051 3289
rect 14874 3273 14983 3278
rect 14874 3261 14915 3273
rect 14807 3239 14915 3261
rect 14949 3244 14983 3273
rect 15017 3255 15051 3278
rect 15085 3255 15100 3289
rect 15017 3244 15100 3255
rect 14949 3239 15100 3244
rect 14807 3227 15100 3239
rect 14807 3193 14840 3227
rect 14874 3217 15100 3227
rect 14874 3205 15051 3217
rect 14874 3200 14983 3205
rect 14874 3193 14915 3200
rect 14807 3166 14915 3193
rect 14949 3171 14983 3200
rect 15017 3183 15051 3205
rect 15085 3183 15100 3217
rect 15017 3171 15100 3183
rect 14949 3166 15100 3171
rect 14807 3159 15100 3166
rect 14807 3125 14840 3159
rect 14874 3145 15100 3159
rect 14874 3132 15051 3145
rect 14874 3127 14983 3132
rect 14874 3125 14915 3127
rect 14807 3093 14915 3125
rect 14949 3098 14983 3127
rect 15017 3111 15051 3132
rect 15085 3111 15100 3145
rect 15017 3098 15100 3111
rect 14949 3093 15100 3098
rect 14807 3091 15100 3093
rect 14807 3057 14840 3091
rect 14874 3073 15100 3091
rect 14874 3059 15051 3073
rect 14874 3057 14983 3059
rect 14807 3054 14983 3057
rect 14807 3023 14915 3054
rect 14807 2989 14840 3023
rect 14874 3020 14915 3023
rect 14949 3025 14983 3054
rect 15017 3039 15051 3059
rect 15085 3039 15100 3073
rect 15017 3025 15100 3039
rect 14949 3020 15100 3025
rect 14874 3001 15100 3020
rect 14874 2989 15051 3001
rect 14807 2986 15051 2989
rect 14807 2981 14983 2986
rect 14807 2955 14915 2981
rect 14807 2921 14840 2955
rect 14874 2947 14915 2955
rect 14949 2952 14983 2981
rect 15017 2967 15051 2986
rect 15085 2967 15100 3001
rect 15017 2952 15100 2967
rect 14949 2947 15100 2952
rect 14874 2929 15100 2947
rect 14874 2921 15051 2929
rect 14807 2913 15051 2921
rect 14807 2908 14983 2913
rect 14807 2887 14915 2908
rect 14807 2853 14840 2887
rect 14874 2874 14915 2887
rect 14949 2879 14983 2908
rect 15017 2895 15051 2913
rect 15085 2895 15100 2929
rect 15017 2879 15100 2895
rect 14949 2874 15100 2879
rect 14874 2857 15100 2874
rect 14874 2853 15051 2857
rect 14807 2840 15051 2853
rect 14807 2835 14983 2840
rect 14807 2819 14915 2835
rect 14807 2785 14840 2819
rect 14874 2801 14915 2819
rect 14949 2806 14983 2835
rect 15017 2823 15051 2840
rect 15085 2823 15100 2857
rect 15017 2806 15100 2823
rect 14949 2801 15100 2806
rect 14874 2785 15100 2801
rect 14807 2767 15051 2785
rect 14807 2762 14983 2767
rect 14807 2751 14915 2762
rect 14807 2717 14840 2751
rect 14874 2728 14915 2751
rect 14949 2733 14983 2762
rect 15017 2751 15051 2767
rect 15085 2751 15100 2785
rect 15017 2733 15100 2751
rect 14949 2728 15100 2733
rect 14874 2717 15100 2728
rect 14807 2713 15100 2717
rect 14807 2694 15051 2713
rect 14807 2689 14983 2694
rect 14807 2683 14915 2689
rect 14807 2649 14840 2683
rect 14874 2655 14915 2683
rect 14949 2660 14983 2689
rect 15017 2679 15051 2694
rect 15085 2679 15100 2713
rect 15017 2660 15100 2679
rect 14949 2655 15100 2660
rect 14874 2649 15100 2655
rect 14807 2641 15100 2649
rect 14807 2621 15051 2641
rect 14807 2616 14983 2621
rect 14807 2615 14915 2616
rect 14807 2581 14840 2615
rect 14874 2582 14915 2615
rect 14949 2587 14983 2616
rect 15017 2607 15051 2621
rect 15085 2607 15100 2641
rect 15017 2587 15100 2607
rect 14949 2582 15100 2587
rect 14874 2581 15100 2582
rect 14807 2569 15100 2581
rect 14807 2548 15051 2569
rect 14807 2547 14983 2548
rect 14807 2513 14840 2547
rect 14874 2543 14983 2547
rect 14874 2513 14915 2543
rect 14807 2509 14915 2513
rect 14949 2514 14983 2543
rect 15017 2535 15051 2548
rect 15085 2535 15100 2569
rect 15017 2514 15100 2535
rect 14949 2509 15100 2514
rect 14807 2497 15100 2509
rect 14807 2479 15051 2497
rect 14807 2445 14840 2479
rect 14874 2475 15051 2479
rect 14874 2470 14983 2475
rect 14874 2445 14915 2470
rect 14807 2436 14915 2445
rect 14949 2441 14983 2470
rect 15017 2463 15051 2475
rect 15085 2463 15100 2497
rect 15017 2441 15100 2463
rect 14949 2436 15100 2441
rect 14807 2425 15100 2436
rect 14807 2411 15051 2425
rect 14807 2377 14840 2411
rect 14874 2402 15051 2411
rect 14874 2397 14983 2402
rect 14874 2377 14915 2397
rect 14807 2363 14915 2377
rect 14949 2368 14983 2397
rect 15017 2391 15051 2402
rect 15085 2391 15100 2425
rect 15017 2368 15100 2391
rect 14949 2363 15100 2368
rect 14807 2353 15100 2363
rect 14807 2343 15051 2353
rect 14807 2309 14840 2343
rect 14874 2329 15051 2343
rect 14874 2324 14983 2329
rect 14874 2309 14915 2324
rect 14807 2290 14915 2309
rect 14949 2295 14983 2324
rect 15017 2319 15051 2329
rect 15085 2319 15100 2353
rect 15017 2295 15100 2319
rect 14949 2290 15100 2295
rect 14807 2280 15100 2290
rect 14807 2275 15051 2280
rect 14807 2241 14840 2275
rect 14874 2256 15051 2275
rect 14874 2251 14983 2256
rect 14874 2241 14915 2251
rect 14807 2217 14915 2241
rect 14949 2222 14983 2251
rect 15017 2246 15051 2256
rect 15085 2246 15100 2280
rect 15017 2222 15100 2246
rect 14949 2217 15100 2222
rect 14807 2207 15100 2217
rect 14807 2173 14840 2207
rect 14874 2183 15051 2207
rect 14874 2178 14983 2183
rect 14874 2173 14915 2178
rect 14807 2144 14915 2173
rect 14949 2149 14983 2178
rect 15017 2173 15051 2183
rect 15085 2173 15100 2207
rect 15017 2149 15100 2173
rect 14949 2144 15100 2149
rect 14807 2139 15100 2144
rect 14807 2105 14840 2139
rect 14874 2134 15100 2139
rect 14874 2110 15051 2134
rect 14874 2105 14983 2110
rect 14807 2071 14915 2105
rect 14949 2076 14983 2105
rect 15017 2100 15051 2110
rect 15085 2100 15100 2134
rect 15017 2076 15100 2100
rect 14949 2071 15100 2076
rect 14807 2037 14840 2071
rect 14874 2061 15100 2071
rect 14874 2037 15051 2061
rect 14807 2032 14983 2037
rect 14807 2003 14915 2032
rect 14807 1969 14840 2003
rect 14874 1998 14915 2003
rect 14949 2003 14983 2032
rect 15017 2027 15051 2037
rect 15085 2027 15100 2061
rect 15017 2003 15100 2027
rect 14949 1998 15100 2003
rect 14874 1988 15100 1998
rect 14874 1969 15051 1988
rect 14807 1964 15051 1969
rect 14807 1959 14983 1964
rect 14807 1935 14915 1959
rect 14807 1901 14840 1935
rect 14874 1925 14915 1935
rect 14949 1930 14983 1959
rect 15017 1954 15051 1964
rect 15085 1954 15100 1988
rect 15017 1930 15100 1954
rect 14949 1925 15100 1930
rect 14874 1915 15100 1925
rect 14874 1901 15051 1915
rect 14807 1891 15051 1901
rect 14807 1886 14983 1891
rect 14807 1867 14915 1886
rect 14807 1833 14840 1867
rect 14874 1852 14915 1867
rect 14949 1857 14983 1886
rect 15017 1881 15051 1891
rect 15085 1881 15100 1915
rect 15017 1857 15100 1881
rect 14949 1852 15100 1857
rect 14874 1842 15100 1852
rect 14874 1833 15051 1842
rect 14807 1818 15051 1833
rect 14807 1813 14983 1818
rect 14807 1799 14915 1813
rect 14807 1765 14840 1799
rect 14874 1779 14915 1799
rect 14949 1784 14983 1813
rect 15017 1808 15051 1818
rect 15085 1808 15100 1842
rect 15017 1784 15100 1808
rect 14949 1779 15100 1784
rect 14874 1769 15100 1779
rect 14874 1765 15051 1769
rect 14807 1745 15051 1765
rect 14807 1740 14983 1745
rect 14807 1731 14915 1740
rect 14807 1697 14840 1731
rect 14874 1706 14915 1731
rect 14949 1711 14983 1740
rect 15017 1735 15051 1745
rect 15085 1735 15100 1769
rect 15017 1711 15100 1735
rect 14949 1706 15100 1711
rect 14874 1697 15100 1706
rect 14807 1696 15100 1697
rect 14807 1672 15051 1696
rect 14807 1667 14983 1672
rect 14807 1663 14915 1667
rect 14807 1629 14840 1663
rect 14874 1633 14915 1663
rect 14949 1638 14983 1667
rect 15017 1662 15051 1672
rect 15085 1662 15100 1696
rect 15017 1638 15100 1662
rect 14949 1633 15100 1638
rect 14874 1629 15100 1633
rect 14807 1623 15100 1629
rect 14807 1599 15051 1623
rect 14807 1595 14983 1599
rect 14807 1561 14840 1595
rect 14874 1594 14983 1595
rect 14874 1561 14915 1594
rect 14807 1560 14915 1561
rect 14949 1565 14983 1594
rect 15017 1589 15051 1599
rect 15085 1589 15100 1623
rect 15017 1565 15100 1589
rect 14949 1560 15100 1565
rect 14807 1550 15100 1560
rect 14807 1527 15051 1550
rect 14807 1493 14840 1527
rect 14874 1526 15051 1527
rect 14874 1521 14983 1526
rect 14874 1493 14915 1521
rect 14807 1487 14915 1493
rect 14949 1492 14983 1521
rect 15017 1516 15051 1526
rect 15085 1516 15100 1550
rect 15017 1492 15100 1516
rect 14949 1487 15100 1492
rect 14807 1477 15100 1487
rect 14807 1459 15051 1477
rect 14807 1425 14840 1459
rect 14874 1453 15051 1459
rect 14874 1448 14983 1453
rect 14874 1425 14915 1448
rect 14807 1414 14915 1425
rect 14949 1419 14983 1448
rect 15017 1443 15051 1453
rect 15085 1443 15100 1477
rect 15017 1419 15100 1443
rect 14949 1414 15100 1419
rect 14807 1404 15100 1414
rect 14807 1391 15051 1404
rect 14807 1357 14840 1391
rect 14874 1380 15051 1391
rect 14874 1375 14983 1380
rect 14874 1357 14915 1375
rect 14807 1341 14915 1357
rect 14949 1346 14983 1375
rect 15017 1370 15051 1380
rect 15085 1370 15100 1404
rect 15017 1346 15100 1370
rect 14949 1341 15100 1346
rect 14807 1331 15100 1341
rect 14807 1323 15051 1331
rect 14807 1289 14840 1323
rect 14874 1307 15051 1323
rect 14874 1302 14983 1307
rect 14874 1289 14915 1302
rect 14807 1268 14915 1289
rect 14949 1273 14983 1302
rect 15017 1297 15051 1307
rect 15085 1297 15100 1331
rect 15017 1273 15100 1297
rect 14949 1268 15100 1273
rect 14807 1258 15100 1268
rect 14807 1255 15051 1258
rect 14807 1221 14840 1255
rect 14874 1234 15051 1255
rect 14874 1229 14983 1234
rect 14874 1221 14915 1229
rect 14807 1195 14915 1221
rect 14949 1200 14983 1229
rect 15017 1224 15051 1234
rect 15085 1224 15100 1258
rect 15017 1200 15100 1224
rect 14949 1195 15100 1200
rect 14807 1187 15100 1195
rect 14807 1153 14840 1187
rect 14874 1185 15100 1187
rect 14874 1161 15051 1185
rect 14874 1156 14983 1161
rect 14874 1153 14915 1156
rect 14807 1122 14915 1153
rect 14949 1127 14983 1156
rect 15017 1151 15051 1161
rect 15085 1151 15100 1185
rect 15017 1127 15100 1151
rect 14949 1122 15100 1127
rect 14807 1119 15100 1122
rect 14807 1085 14840 1119
rect 14874 1112 15100 1119
rect 14874 1088 15051 1112
rect 14874 1085 14983 1088
rect 14807 1083 14983 1085
rect 14807 1051 14915 1083
rect 14807 1017 14840 1051
rect 14874 1049 14915 1051
rect 14949 1054 14983 1083
rect 15017 1078 15051 1088
rect 15085 1078 15100 1112
rect 15017 1054 15100 1078
rect 14949 1049 15100 1054
rect 14874 1039 15100 1049
rect 14874 1017 15051 1039
rect 14807 1015 15051 1017
rect 14807 1010 14983 1015
rect 14807 983 14915 1010
rect 14807 949 14840 983
rect 14874 976 14915 983
rect 14949 981 14983 1010
rect 15017 1005 15051 1015
rect 15085 1005 15100 1039
rect 15017 981 15100 1005
rect 14949 976 15100 981
rect 14874 966 15100 976
rect 14874 949 15051 966
rect 14807 942 15051 949
rect 14807 937 14983 942
rect 14807 915 14915 937
rect 14807 881 14840 915
rect 14874 903 14915 915
rect 14949 908 14983 937
rect 15017 932 15051 942
rect 15085 932 15100 966
rect 15017 908 15100 932
rect 14949 903 15100 908
rect 14874 893 15100 903
rect 14874 881 15051 893
rect 14807 869 15051 881
rect 14807 864 14983 869
rect 14807 847 14915 864
rect 14807 813 14840 847
rect 14874 830 14915 847
rect 14949 835 14983 864
rect 15017 859 15051 869
rect 15085 859 15100 893
rect 15017 835 15100 859
rect 14949 830 15100 835
rect 14874 820 15100 830
rect 14874 813 15051 820
rect 14807 796 15051 813
rect 14807 791 14983 796
rect 14807 779 14915 791
rect 14807 745 14840 779
rect 14874 757 14915 779
rect 14949 762 14983 791
rect 15017 786 15051 796
rect 15085 786 15100 820
rect 15017 762 15100 786
rect 14949 757 15100 762
rect 14874 747 15100 757
rect 14874 745 15051 747
rect 14807 723 15051 745
rect 14807 718 14983 723
rect 14807 711 14915 718
rect 14807 677 14840 711
rect 14874 684 14915 711
rect 14949 689 14983 718
rect 15017 713 15051 723
rect 15085 713 15100 747
rect 15017 689 15100 713
rect 14949 684 15100 689
rect 14874 677 15100 684
rect 14807 674 15100 677
rect 36 643 329 648
rect 36 610 262 643
rect 36 576 51 610
rect 85 576 119 610
rect 153 576 187 610
rect 221 609 262 610
rect 296 609 329 643
rect 221 576 329 609
rect 36 575 329 576
rect 36 541 262 575
rect 296 541 329 575
rect 36 538 329 541
rect 36 504 51 538
rect 85 504 119 538
rect 153 504 187 538
rect 221 514 329 538
rect 14807 650 15051 674
rect 14807 645 14983 650
rect 14807 643 14915 645
rect 14807 609 14840 643
rect 14874 611 14915 643
rect 14949 616 14983 645
rect 15017 640 15051 650
rect 15085 640 15100 674
rect 15017 616 15100 640
rect 14949 611 15100 616
rect 14874 609 15100 611
rect 14807 601 15100 609
rect 14807 577 15051 601
rect 14807 575 14983 577
rect 14807 541 14840 575
rect 14874 572 14983 575
rect 14874 541 14915 572
rect 14807 538 14915 541
rect 14949 543 14983 572
rect 15017 567 15051 577
rect 15085 567 15100 601
rect 15017 543 15100 567
rect 14949 538 15100 543
rect 14807 528 15100 538
rect 14807 514 15051 528
rect 221 504 15051 514
rect 36 499 14983 504
rect 36 466 302 499
rect 36 432 51 466
rect 85 432 119 466
rect 153 432 187 466
rect 221 465 302 466
rect 336 465 375 499
rect 409 465 448 499
rect 482 465 521 499
rect 555 465 594 499
rect 628 465 667 499
rect 701 465 740 499
rect 774 465 813 499
rect 847 465 886 499
rect 920 465 959 499
rect 993 465 1032 499
rect 1066 465 1105 499
rect 1139 465 1178 499
rect 1212 465 1251 499
rect 1285 465 1324 499
rect 1358 465 1397 499
rect 1431 465 1470 499
rect 1504 465 1543 499
rect 1577 465 1616 499
rect 1650 465 1689 499
rect 1723 465 1762 499
rect 1796 465 1835 499
rect 1869 465 1908 499
rect 1942 465 1981 499
rect 2015 465 2054 499
rect 2088 465 2127 499
rect 2161 465 2200 499
rect 2234 465 2273 499
rect 2307 465 2346 499
rect 2380 465 2419 499
rect 2453 465 2492 499
rect 2526 465 2565 499
rect 2599 465 2638 499
rect 2672 465 2711 499
rect 2745 465 2784 499
rect 2818 465 2857 499
rect 2891 465 2930 499
rect 2964 465 3003 499
rect 3037 465 3076 499
rect 3110 465 3149 499
rect 3183 465 3222 499
rect 3256 465 3295 499
rect 3329 465 3368 499
rect 3402 465 3441 499
rect 3475 465 3514 499
rect 3548 465 3587 499
rect 3621 465 3660 499
rect 3694 465 3733 499
rect 3767 465 3806 499
rect 3840 465 3879 499
rect 3913 465 3952 499
rect 3986 465 4025 499
rect 4059 465 4098 499
rect 4132 465 4171 499
rect 4205 465 4244 499
rect 4278 465 4317 499
rect 4351 465 4390 499
rect 4424 465 4463 499
rect 4497 465 4536 499
rect 4570 465 4609 499
rect 4643 465 4682 499
rect 4716 465 4755 499
rect 4789 465 4828 499
rect 4862 465 4901 499
rect 4935 465 4974 499
rect 5008 465 5047 499
rect 5081 465 5120 499
rect 5154 465 5193 499
rect 5227 465 5266 499
rect 5300 465 5339 499
rect 5373 465 5411 499
rect 5445 465 5483 499
rect 5517 465 5555 499
rect 5589 465 5627 499
rect 5661 465 5699 499
rect 5733 465 5771 499
rect 5805 465 5843 499
rect 5877 465 5915 499
rect 5949 465 5987 499
rect 6021 465 6059 499
rect 6093 465 6131 499
rect 6165 465 6203 499
rect 6237 465 6275 499
rect 6309 465 6347 499
rect 6381 465 6419 499
rect 6453 465 6491 499
rect 6525 465 6563 499
rect 6597 465 6635 499
rect 6669 465 6707 499
rect 6741 465 6779 499
rect 6813 465 6851 499
rect 6885 465 6923 499
rect 6957 465 6995 499
rect 7029 465 7067 499
rect 7101 465 7139 499
rect 7173 465 7211 499
rect 7245 465 7283 499
rect 7317 465 7355 499
rect 7389 465 7427 499
rect 7461 465 7499 499
rect 7533 465 7571 499
rect 7605 465 7643 499
rect 7677 465 7715 499
rect 7749 465 7787 499
rect 7821 465 7859 499
rect 7893 465 7931 499
rect 7965 465 8003 499
rect 8037 465 8075 499
rect 8109 465 8147 499
rect 8181 465 8219 499
rect 8253 465 8291 499
rect 8325 465 8363 499
rect 8397 465 8435 499
rect 8469 465 8507 499
rect 8541 465 8579 499
rect 8613 465 8651 499
rect 8685 465 8723 499
rect 8757 465 8795 499
rect 8829 465 8867 499
rect 8901 465 8939 499
rect 8973 465 9011 499
rect 9045 465 9083 499
rect 9117 465 9155 499
rect 9189 465 9227 499
rect 9261 465 9299 499
rect 9333 465 9371 499
rect 9405 465 9443 499
rect 9477 465 9515 499
rect 9549 465 9587 499
rect 9621 465 9659 499
rect 9693 465 9731 499
rect 9765 465 9803 499
rect 9837 465 9875 499
rect 9909 465 9947 499
rect 9981 465 10019 499
rect 10053 465 10091 499
rect 10125 465 10163 499
rect 10197 465 10235 499
rect 10269 465 10307 499
rect 10341 465 10379 499
rect 10413 465 10451 499
rect 10485 465 10523 499
rect 10557 465 10595 499
rect 10629 465 10667 499
rect 10701 465 10739 499
rect 10773 465 10811 499
rect 10845 465 10883 499
rect 10917 465 10955 499
rect 10989 465 11027 499
rect 11061 465 11099 499
rect 11133 465 11171 499
rect 11205 465 11243 499
rect 11277 465 11315 499
rect 11349 465 11387 499
rect 11421 465 11459 499
rect 11493 465 11531 499
rect 11565 465 11603 499
rect 11637 465 11675 499
rect 11709 465 11747 499
rect 11781 465 11819 499
rect 11853 465 11891 499
rect 11925 465 11963 499
rect 11997 465 12035 499
rect 12069 465 12107 499
rect 12141 465 12179 499
rect 12213 465 12251 499
rect 12285 465 12323 499
rect 12357 465 12395 499
rect 12429 465 12467 499
rect 12501 465 12539 499
rect 12573 465 12611 499
rect 12645 465 12683 499
rect 12717 465 12755 499
rect 12789 465 12827 499
rect 12861 465 12899 499
rect 12933 465 12971 499
rect 13005 465 13043 499
rect 13077 465 13115 499
rect 13149 465 13187 499
rect 13221 465 13259 499
rect 13293 465 13331 499
rect 13365 465 13403 499
rect 13437 465 13475 499
rect 13509 465 13547 499
rect 13581 465 13619 499
rect 13653 465 13691 499
rect 13725 465 13763 499
rect 13797 465 13835 499
rect 13869 465 13907 499
rect 13941 465 13979 499
rect 14013 465 14051 499
rect 14085 465 14123 499
rect 14157 465 14195 499
rect 14229 465 14267 499
rect 14301 465 14339 499
rect 14373 465 14411 499
rect 14445 465 14483 499
rect 14517 465 14555 499
rect 14589 465 14627 499
rect 14661 465 14699 499
rect 14733 465 14771 499
rect 14805 465 14843 499
rect 14877 465 14915 499
rect 14949 470 14983 499
rect 15017 494 15051 504
rect 15085 494 15100 528
rect 15017 470 15100 494
rect 14949 465 15100 470
rect 221 455 15100 465
rect 221 432 15051 455
rect 36 431 15051 432
rect 36 397 302 431
rect 336 397 375 431
rect 409 397 448 431
rect 482 397 521 431
rect 555 397 594 431
rect 628 397 667 431
rect 701 397 740 431
rect 774 397 813 431
rect 847 397 886 431
rect 920 397 959 431
rect 993 397 1032 431
rect 1066 397 1105 431
rect 1139 397 1178 431
rect 1212 397 1251 431
rect 1285 397 1324 431
rect 1358 397 1397 431
rect 1431 397 1470 431
rect 1504 397 1543 431
rect 1577 397 1616 431
rect 1650 397 1689 431
rect 1723 397 1762 431
rect 1796 397 1835 431
rect 1869 397 1908 431
rect 1942 397 1981 431
rect 2015 397 2054 431
rect 2088 397 2127 431
rect 2161 397 2200 431
rect 2234 397 2273 431
rect 2307 397 2346 431
rect 2380 397 2419 431
rect 2453 397 2492 431
rect 2526 397 2565 431
rect 2599 397 2638 431
rect 2672 397 2711 431
rect 2745 397 2784 431
rect 2818 397 2857 431
rect 2891 397 2930 431
rect 2964 397 3003 431
rect 3037 397 3076 431
rect 3110 397 3149 431
rect 3183 397 3222 431
rect 3256 397 3295 431
rect 3329 397 3368 431
rect 3402 397 3441 431
rect 3475 397 3514 431
rect 3548 397 3587 431
rect 3621 397 3660 431
rect 3694 397 3733 431
rect 3767 397 3806 431
rect 3840 397 3879 431
rect 3913 397 3952 431
rect 3986 397 4025 431
rect 4059 397 4098 431
rect 4132 397 4171 431
rect 4205 397 4244 431
rect 4278 397 4317 431
rect 4351 397 4390 431
rect 4424 397 4463 431
rect 4497 397 4536 431
rect 4570 397 4609 431
rect 4643 397 4682 431
rect 4716 397 4755 431
rect 4789 397 4828 431
rect 4862 397 4901 431
rect 4935 397 4974 431
rect 5008 397 5047 431
rect 5081 397 5119 431
rect 5153 397 5191 431
rect 5225 397 5263 431
rect 5297 397 5335 431
rect 5369 397 5407 431
rect 5441 397 5479 431
rect 5513 397 5551 431
rect 5585 397 5623 431
rect 5657 397 5695 431
rect 5729 397 5767 431
rect 5801 397 5839 431
rect 5873 397 5911 431
rect 5945 397 5983 431
rect 6017 397 6055 431
rect 6089 397 6127 431
rect 6161 397 6199 431
rect 6233 397 6271 431
rect 6305 397 6343 431
rect 6377 397 6415 431
rect 6449 397 6487 431
rect 6521 397 6559 431
rect 6593 397 6631 431
rect 6665 397 6703 431
rect 6737 397 6775 431
rect 6809 397 6847 431
rect 6881 397 6919 431
rect 6953 397 6991 431
rect 7025 397 7063 431
rect 7097 397 7135 431
rect 7169 397 7207 431
rect 7241 397 7279 431
rect 7313 397 7351 431
rect 7385 397 7423 431
rect 7457 397 7495 431
rect 7529 397 7567 431
rect 7601 397 7639 431
rect 7673 397 7711 431
rect 7745 397 7783 431
rect 7817 397 7855 431
rect 7889 397 7927 431
rect 7961 397 7999 431
rect 8033 397 8071 431
rect 8105 397 8143 431
rect 8177 397 8215 431
rect 8249 397 8287 431
rect 8321 397 8359 431
rect 8393 397 8431 431
rect 8465 397 8503 431
rect 8537 397 8575 431
rect 8609 397 8647 431
rect 8681 397 8719 431
rect 8753 397 8791 431
rect 8825 397 8863 431
rect 8897 397 8935 431
rect 8969 397 9007 431
rect 9041 397 9079 431
rect 9113 397 9151 431
rect 9185 397 9223 431
rect 9257 397 9295 431
rect 9329 397 9367 431
rect 9401 397 9439 431
rect 9473 397 9511 431
rect 9545 397 9583 431
rect 9617 397 9655 431
rect 9689 397 9727 431
rect 9761 397 9799 431
rect 9833 397 9871 431
rect 9905 397 9943 431
rect 9977 397 10015 431
rect 10049 397 10087 431
rect 10121 397 10159 431
rect 10193 397 10231 431
rect 10265 397 10303 431
rect 10337 397 10375 431
rect 10409 397 10447 431
rect 10481 397 10519 431
rect 10553 397 10591 431
rect 10625 397 10663 431
rect 10697 397 10735 431
rect 10769 397 10807 431
rect 10841 397 10879 431
rect 10913 397 10951 431
rect 10985 397 11023 431
rect 11057 397 11095 431
rect 11129 397 11167 431
rect 11201 397 11239 431
rect 11273 397 11311 431
rect 11345 397 11383 431
rect 11417 397 11455 431
rect 11489 397 11527 431
rect 11561 397 11599 431
rect 11633 397 11671 431
rect 11705 397 11743 431
rect 11777 397 11815 431
rect 11849 397 11887 431
rect 11921 397 11959 431
rect 11993 397 12031 431
rect 12065 397 12103 431
rect 12137 397 12175 431
rect 12209 397 12247 431
rect 12281 397 12319 431
rect 12353 397 12391 431
rect 12425 397 12463 431
rect 12497 397 12535 431
rect 12569 397 12607 431
rect 12641 397 12679 431
rect 12713 397 12751 431
rect 12785 397 12823 431
rect 12857 397 12895 431
rect 12929 397 12967 431
rect 13001 397 13039 431
rect 13073 397 13111 431
rect 13145 397 13183 431
rect 13217 397 13255 431
rect 13289 397 13327 431
rect 13361 397 13399 431
rect 13433 397 13471 431
rect 13505 397 13543 431
rect 13577 397 13615 431
rect 13649 397 13687 431
rect 13721 397 13759 431
rect 13793 397 13831 431
rect 13865 397 13903 431
rect 13937 397 13975 431
rect 14009 397 14047 431
rect 14081 397 14119 431
rect 14153 397 14191 431
rect 14225 397 14263 431
rect 14297 397 14335 431
rect 14369 397 14407 431
rect 14441 397 14479 431
rect 14513 397 14551 431
rect 14585 397 14623 431
rect 14657 397 14695 431
rect 14729 397 14767 431
rect 14801 397 14839 431
rect 14873 397 14911 431
rect 14945 397 14983 431
rect 15017 421 15051 431
rect 15085 421 15100 455
rect 15017 397 15100 421
rect 36 394 15100 397
rect 36 360 51 394
rect 85 360 119 394
rect 153 360 187 394
rect 221 382 15100 394
rect 221 363 15051 382
rect 221 360 302 363
rect 36 329 302 360
rect 336 329 375 363
rect 409 329 448 363
rect 482 329 521 363
rect 555 329 594 363
rect 628 329 667 363
rect 701 329 740 363
rect 774 329 813 363
rect 847 329 886 363
rect 920 329 959 363
rect 993 329 1032 363
rect 1066 329 1105 363
rect 1139 329 1178 363
rect 1212 329 1251 363
rect 1285 329 1324 363
rect 1358 329 1397 363
rect 1431 329 1470 363
rect 1504 329 1543 363
rect 1577 329 1616 363
rect 1650 329 1689 363
rect 1723 329 1762 363
rect 1796 329 1835 363
rect 1869 329 1908 363
rect 1942 329 1981 363
rect 2015 329 2054 363
rect 2088 329 2127 363
rect 2161 329 2200 363
rect 2234 329 2273 363
rect 2307 329 2346 363
rect 2380 329 2419 363
rect 2453 329 2492 363
rect 2526 329 2565 363
rect 2599 329 2638 363
rect 2672 329 2711 363
rect 2745 329 2784 363
rect 2818 329 2857 363
rect 2891 329 2930 363
rect 2964 329 3003 363
rect 3037 329 3076 363
rect 3110 329 3149 363
rect 3183 329 3222 363
rect 3256 329 3295 363
rect 3329 329 3368 363
rect 3402 329 3440 363
rect 3474 329 3512 363
rect 3546 329 3584 363
rect 3618 329 3656 363
rect 3690 329 3728 363
rect 3762 329 3800 363
rect 3834 329 3872 363
rect 3906 329 3944 363
rect 3978 329 4016 363
rect 4050 329 4088 363
rect 4122 329 4160 363
rect 4194 329 4232 363
rect 4266 329 4304 363
rect 4338 329 4376 363
rect 4410 329 4448 363
rect 4482 329 4520 363
rect 4554 329 4592 363
rect 4626 329 4664 363
rect 4698 329 4736 363
rect 4770 329 4808 363
rect 4842 329 4880 363
rect 4914 329 4952 363
rect 4986 329 5024 363
rect 5058 329 5096 363
rect 5130 329 5168 363
rect 5202 329 5240 363
rect 5274 329 5312 363
rect 5346 329 5384 363
rect 5418 329 5456 363
rect 5490 329 5528 363
rect 5562 329 5600 363
rect 5634 329 5672 363
rect 5706 329 5744 363
rect 5778 329 5816 363
rect 5850 329 5888 363
rect 5922 329 5960 363
rect 5994 329 6032 363
rect 6066 329 6104 363
rect 6138 329 6176 363
rect 6210 329 6248 363
rect 6282 329 6320 363
rect 6354 329 6392 363
rect 6426 329 6464 363
rect 6498 329 6536 363
rect 6570 329 6608 363
rect 6642 329 6680 363
rect 6714 329 6752 363
rect 6786 329 6824 363
rect 6858 329 6896 363
rect 6930 329 6968 363
rect 7002 329 7040 363
rect 7074 329 7112 363
rect 7146 329 7184 363
rect 7218 329 7256 363
rect 7290 329 7328 363
rect 7362 329 7400 363
rect 7434 329 7472 363
rect 7506 329 7544 363
rect 7578 329 7616 363
rect 7650 329 7688 363
rect 7722 329 7760 363
rect 7794 329 7832 363
rect 7866 329 7904 363
rect 7938 329 7976 363
rect 8010 329 8048 363
rect 8082 329 8120 363
rect 8154 329 8192 363
rect 8226 329 8264 363
rect 8298 329 8336 363
rect 8370 329 8408 363
rect 8442 329 8480 363
rect 8514 329 8552 363
rect 8586 329 8624 363
rect 8658 329 8696 363
rect 8730 329 8768 363
rect 8802 329 8840 363
rect 8874 329 8912 363
rect 8946 329 8984 363
rect 9018 329 9056 363
rect 9090 329 9128 363
rect 9162 329 9200 363
rect 9234 329 9272 363
rect 9306 329 9344 363
rect 9378 329 9416 363
rect 9450 329 9488 363
rect 9522 329 9560 363
rect 9594 329 9632 363
rect 9666 329 9704 363
rect 9738 329 9776 363
rect 9810 329 9848 363
rect 9882 329 9920 363
rect 9954 329 9992 363
rect 10026 329 10064 363
rect 10098 329 10136 363
rect 10170 329 10208 363
rect 10242 329 10280 363
rect 10314 329 10352 363
rect 10386 329 10424 363
rect 10458 329 10496 363
rect 10530 329 10568 363
rect 10602 329 10640 363
rect 10674 329 10712 363
rect 10746 329 10784 363
rect 10818 329 10856 363
rect 10890 329 10928 363
rect 10962 329 11000 363
rect 11034 329 11072 363
rect 11106 329 11144 363
rect 11178 329 11216 363
rect 11250 329 11288 363
rect 11322 329 11360 363
rect 11394 329 11432 363
rect 11466 329 11504 363
rect 11538 329 11576 363
rect 11610 329 11648 363
rect 11682 329 11720 363
rect 11754 329 11792 363
rect 11826 329 11864 363
rect 11898 329 11936 363
rect 11970 329 12008 363
rect 12042 329 12080 363
rect 12114 329 12152 363
rect 12186 329 12224 363
rect 12258 329 12296 363
rect 12330 329 12368 363
rect 12402 329 12440 363
rect 12474 329 12512 363
rect 12546 329 12584 363
rect 12618 329 12656 363
rect 12690 329 12728 363
rect 12762 329 12800 363
rect 12834 329 12872 363
rect 12906 329 12944 363
rect 12978 329 13016 363
rect 13050 329 13088 363
rect 13122 329 13160 363
rect 13194 329 13232 363
rect 13266 329 13304 363
rect 13338 329 13376 363
rect 13410 329 13448 363
rect 13482 329 13520 363
rect 13554 329 13592 363
rect 13626 329 13664 363
rect 13698 329 13736 363
rect 13770 329 13808 363
rect 13842 329 13880 363
rect 13914 329 13952 363
rect 13986 329 14024 363
rect 14058 329 14096 363
rect 14130 329 14168 363
rect 14202 329 14240 363
rect 14274 329 14312 363
rect 14346 329 14384 363
rect 14418 329 14456 363
rect 14490 329 14528 363
rect 14562 329 14600 363
rect 14634 329 14672 363
rect 14706 329 14744 363
rect 14778 329 14816 363
rect 14850 329 14888 363
rect 14922 329 14960 363
rect 14994 348 15051 363
rect 15085 348 15100 382
rect 14994 329 15100 348
rect 36 314 15100 329
<< mvnsubdiff >>
rect 482 4638 14653 4653
rect 482 4619 584 4638
rect 482 4585 497 4619
rect 531 4585 584 4619
rect 482 4570 584 4585
rect 10410 4604 10445 4638
rect 10479 4604 10514 4638
rect 10548 4604 10583 4638
rect 10617 4604 10652 4638
rect 10686 4604 10721 4638
rect 10755 4604 10790 4638
rect 10824 4604 10859 4638
rect 10893 4604 10928 4638
rect 10962 4604 10997 4638
rect 11031 4604 11066 4638
rect 11100 4604 11135 4638
rect 11169 4604 11204 4638
rect 11238 4604 11273 4638
rect 11307 4604 11342 4638
rect 11376 4604 11411 4638
rect 11445 4604 11480 4638
rect 11514 4604 11549 4638
rect 11583 4604 11618 4638
rect 11652 4604 11687 4638
rect 11721 4604 11756 4638
rect 11790 4604 11825 4638
rect 11859 4604 11894 4638
rect 11928 4604 11963 4638
rect 11997 4604 12032 4638
rect 12066 4604 12101 4638
rect 12135 4604 12170 4638
rect 12204 4604 12239 4638
rect 12273 4604 12308 4638
rect 12342 4604 12377 4638
rect 12411 4604 12446 4638
rect 12480 4604 12515 4638
rect 12549 4604 12584 4638
rect 12618 4604 12653 4638
rect 12687 4604 12722 4638
rect 12756 4604 12791 4638
rect 12825 4604 12860 4638
rect 12894 4604 12929 4638
rect 12963 4604 12998 4638
rect 13032 4604 13067 4638
rect 13101 4604 13136 4638
rect 13170 4604 13205 4638
rect 13239 4604 13274 4638
rect 13308 4604 13343 4638
rect 13377 4604 13412 4638
rect 13446 4604 13481 4638
rect 13515 4604 13550 4638
rect 13584 4604 13619 4638
rect 13653 4604 13688 4638
rect 13722 4604 13757 4638
rect 13791 4604 13826 4638
rect 13860 4604 13895 4638
rect 13929 4604 13964 4638
rect 13998 4604 14033 4638
rect 14067 4604 14102 4638
rect 14136 4604 14171 4638
rect 14205 4604 14240 4638
rect 14274 4604 14309 4638
rect 14343 4604 14378 4638
rect 14412 4604 14447 4638
rect 14481 4604 14516 4638
rect 14550 4604 14585 4638
rect 14619 4604 14653 4638
rect 10410 4570 14653 4604
rect 482 4549 565 4570
rect 482 4515 497 4549
rect 531 4536 565 4549
rect 12363 4536 12397 4570
rect 12431 4536 12466 4570
rect 12500 4536 12535 4570
rect 12569 4536 12604 4570
rect 12638 4536 12673 4570
rect 12707 4536 12742 4570
rect 12776 4536 12811 4570
rect 12845 4536 12880 4570
rect 12914 4536 12949 4570
rect 12983 4536 13018 4570
rect 13052 4536 13087 4570
rect 13121 4536 13156 4570
rect 13190 4536 13225 4570
rect 13259 4536 13294 4570
rect 13328 4536 13363 4570
rect 13397 4536 13432 4570
rect 13466 4536 13501 4570
rect 13535 4536 13570 4570
rect 13604 4536 13639 4570
rect 13673 4536 13708 4570
rect 13742 4536 13777 4570
rect 13811 4536 13846 4570
rect 13880 4536 13915 4570
rect 13949 4536 13984 4570
rect 14018 4536 14053 4570
rect 14087 4536 14122 4570
rect 14156 4536 14191 4570
rect 14225 4536 14260 4570
rect 14294 4536 14329 4570
rect 14363 4536 14398 4570
rect 14432 4536 14467 4570
rect 14501 4536 14536 4570
rect 14570 4551 14653 4570
rect 531 4515 633 4536
rect 482 4498 633 4515
rect 482 4479 565 4498
rect 482 4445 497 4479
rect 531 4464 565 4479
rect 599 4468 633 4498
rect 12363 4502 14536 4536
rect 12363 4468 12398 4502
rect 12432 4468 12467 4502
rect 12501 4468 12536 4502
rect 12570 4468 12605 4502
rect 12639 4468 12674 4502
rect 12708 4468 12743 4502
rect 12777 4468 12812 4502
rect 12846 4468 12881 4502
rect 12915 4468 12950 4502
rect 12984 4468 13019 4502
rect 13053 4468 13088 4502
rect 13122 4468 13157 4502
rect 13191 4468 13226 4502
rect 13260 4468 13295 4502
rect 13329 4468 13364 4502
rect 13398 4468 13433 4502
rect 13467 4468 13502 4502
rect 13536 4468 13571 4502
rect 13605 4468 13640 4502
rect 13674 4468 13709 4502
rect 13743 4468 13778 4502
rect 13812 4468 13847 4502
rect 13881 4468 13916 4502
rect 13950 4468 13985 4502
rect 14019 4468 14054 4502
rect 14088 4468 14123 4502
rect 14157 4468 14192 4502
rect 14226 4468 14261 4502
rect 14295 4468 14330 4502
rect 14364 4468 14399 4502
rect 14433 4468 14468 4502
rect 599 4464 14468 4468
rect 531 4453 14468 4464
rect 531 4445 682 4453
rect 482 4429 682 4445
rect 482 4426 633 4429
rect 482 4409 565 4426
rect 482 4375 497 4409
rect 531 4392 565 4409
rect 599 4395 633 4426
rect 667 4395 682 4429
rect 599 4392 682 4395
rect 531 4375 682 4392
rect 482 4356 682 4375
rect 482 4354 633 4356
rect 482 4339 565 4354
rect 482 4305 497 4339
rect 531 4320 565 4339
rect 599 4322 633 4354
rect 667 4322 682 4356
rect 599 4320 682 4322
rect 531 4305 682 4320
rect 482 4283 682 4305
rect 482 4282 633 4283
rect 482 4269 565 4282
rect 482 4235 497 4269
rect 531 4248 565 4269
rect 599 4249 633 4282
rect 667 4249 682 4283
rect 599 4248 682 4249
rect 531 4235 682 4248
rect 482 4211 682 4235
rect 482 4210 633 4211
rect 482 4199 565 4210
rect 482 4165 497 4199
rect 531 4176 565 4199
rect 599 4177 633 4210
rect 667 4177 682 4211
rect 599 4176 682 4177
rect 531 4165 682 4176
rect 482 4152 682 4165
rect 14453 4152 14468 4453
rect 482 4139 708 4152
rect 482 4138 633 4139
rect 482 4129 565 4138
rect 482 4095 497 4129
rect 531 4104 565 4129
rect 599 4105 633 4138
rect 667 4105 708 4139
rect 599 4104 708 4105
rect 531 4095 708 4104
rect 482 4067 708 4095
rect 482 4066 633 4067
rect 482 4059 565 4066
rect 482 4025 497 4059
rect 531 4032 565 4059
rect 599 4033 633 4066
rect 667 4033 708 4067
rect 599 4032 708 4033
rect 531 4025 708 4032
rect 482 3995 708 4025
rect 482 3994 633 3995
rect 482 3989 565 3994
rect 482 3955 497 3989
rect 531 3960 565 3989
rect 599 3961 633 3994
rect 667 3961 708 3995
rect 599 3960 708 3961
rect 531 3955 708 3960
rect 482 3923 708 3955
rect 482 3922 633 3923
rect 482 3920 565 3922
rect 482 3886 497 3920
rect 531 3888 565 3920
rect 599 3889 633 3922
rect 667 3889 708 3923
rect 599 3888 708 3889
rect 531 3886 708 3888
rect 482 3851 708 3886
rect 482 3817 497 3851
rect 531 3817 565 3851
rect 599 3817 633 3851
rect 667 3817 708 3851
rect 482 3749 708 3817
rect 482 3715 497 3749
rect 531 3715 565 3749
rect 599 3715 633 3749
rect 667 3715 708 3749
rect 482 3680 708 3715
rect 482 3646 497 3680
rect 531 3646 565 3680
rect 599 3646 633 3680
rect 667 3646 708 3680
rect 482 3611 708 3646
rect 482 3577 497 3611
rect 531 3577 565 3611
rect 599 3577 633 3611
rect 667 3577 708 3611
rect 482 3542 708 3577
rect 482 3508 497 3542
rect 531 3508 565 3542
rect 599 3508 633 3542
rect 667 3508 708 3542
rect 482 3473 708 3508
rect 482 3439 497 3473
rect 531 3439 565 3473
rect 599 3439 633 3473
rect 667 3439 708 3473
rect 482 3404 708 3439
rect 482 3370 497 3404
rect 531 3370 565 3404
rect 599 3370 633 3404
rect 667 3370 708 3404
rect 482 3335 708 3370
rect 482 3301 497 3335
rect 531 3301 565 3335
rect 599 3301 633 3335
rect 667 3301 708 3335
rect 482 3266 708 3301
rect 482 3232 497 3266
rect 531 3232 565 3266
rect 599 3232 633 3266
rect 667 3232 708 3266
rect 482 3197 708 3232
rect 482 3163 497 3197
rect 531 3163 565 3197
rect 599 3163 633 3197
rect 667 3163 708 3197
rect 482 3152 708 3163
rect 1582 4082 1722 4152
rect 1582 4048 1635 4082
rect 1669 4048 1722 4082
rect 1582 4014 1722 4048
rect 1582 3980 1635 4014
rect 1669 3980 1722 4014
rect 1582 3946 1722 3980
rect 1582 3912 1635 3946
rect 1669 3912 1722 3946
rect 1582 3878 1722 3912
rect 1582 3844 1635 3878
rect 1669 3844 1722 3878
rect 1582 3810 1722 3844
rect 1582 3776 1635 3810
rect 1669 3776 1722 3810
rect 1582 3742 1722 3776
rect 1582 3708 1635 3742
rect 1669 3708 1722 3742
rect 1582 3674 1722 3708
rect 1582 3640 1635 3674
rect 1669 3640 1722 3674
rect 1582 3606 1722 3640
rect 1582 3572 1635 3606
rect 1669 3572 1722 3606
rect 1582 3538 1722 3572
rect 1582 3504 1635 3538
rect 1669 3504 1722 3538
rect 1582 3470 1722 3504
rect 1582 3436 1635 3470
rect 1669 3436 1722 3470
rect 1582 3402 1722 3436
rect 1582 3368 1635 3402
rect 1669 3368 1722 3402
rect 1582 3334 1722 3368
rect 1582 3300 1635 3334
rect 1669 3300 1722 3334
rect 1582 3266 1722 3300
rect 1582 3232 1635 3266
rect 1669 3232 1722 3266
rect 1582 3198 1722 3232
rect 1582 3164 1635 3198
rect 1669 3164 1722 3198
rect 1582 3152 1722 3164
rect 2574 4082 2714 4152
rect 2574 4048 2627 4082
rect 2661 4048 2714 4082
rect 2574 4014 2714 4048
rect 2574 3980 2627 4014
rect 2661 3980 2714 4014
rect 2574 3946 2714 3980
rect 2574 3912 2627 3946
rect 2661 3912 2714 3946
rect 2574 3878 2714 3912
rect 2574 3844 2627 3878
rect 2661 3844 2714 3878
rect 2574 3810 2714 3844
rect 2574 3776 2627 3810
rect 2661 3776 2714 3810
rect 2574 3742 2714 3776
rect 2574 3708 2627 3742
rect 2661 3708 2714 3742
rect 2574 3674 2714 3708
rect 2574 3640 2627 3674
rect 2661 3640 2714 3674
rect 2574 3606 2714 3640
rect 2574 3572 2627 3606
rect 2661 3572 2714 3606
rect 2574 3538 2714 3572
rect 2574 3504 2627 3538
rect 2661 3504 2714 3538
rect 2574 3470 2714 3504
rect 2574 3436 2627 3470
rect 2661 3436 2714 3470
rect 2574 3402 2714 3436
rect 2574 3368 2627 3402
rect 2661 3368 2714 3402
rect 2574 3334 2714 3368
rect 2574 3300 2627 3334
rect 2661 3300 2714 3334
rect 2574 3266 2714 3300
rect 2574 3232 2627 3266
rect 2661 3232 2714 3266
rect 2574 3198 2714 3232
rect 2574 3164 2627 3198
rect 2661 3164 2714 3198
rect 2574 3152 2714 3164
rect 3566 4082 3706 4152
rect 3566 4048 3619 4082
rect 3653 4048 3706 4082
rect 3566 4014 3706 4048
rect 3566 3980 3619 4014
rect 3653 3980 3706 4014
rect 3566 3946 3706 3980
rect 3566 3912 3619 3946
rect 3653 3912 3706 3946
rect 3566 3878 3706 3912
rect 3566 3844 3619 3878
rect 3653 3844 3706 3878
rect 3566 3810 3706 3844
rect 3566 3776 3619 3810
rect 3653 3776 3706 3810
rect 3566 3742 3706 3776
rect 3566 3708 3619 3742
rect 3653 3708 3706 3742
rect 3566 3674 3706 3708
rect 3566 3640 3619 3674
rect 3653 3640 3706 3674
rect 3566 3606 3706 3640
rect 3566 3572 3619 3606
rect 3653 3572 3706 3606
rect 3566 3538 3706 3572
rect 3566 3504 3619 3538
rect 3653 3504 3706 3538
rect 3566 3470 3706 3504
rect 3566 3436 3619 3470
rect 3653 3436 3706 3470
rect 3566 3402 3706 3436
rect 3566 3368 3619 3402
rect 3653 3368 3706 3402
rect 3566 3334 3706 3368
rect 3566 3300 3619 3334
rect 3653 3300 3706 3334
rect 3566 3266 3706 3300
rect 3566 3232 3619 3266
rect 3653 3232 3706 3266
rect 3566 3198 3706 3232
rect 3566 3164 3619 3198
rect 3653 3164 3706 3198
rect 3566 3152 3706 3164
rect 4558 4082 4698 4152
rect 4558 4048 4611 4082
rect 4645 4048 4698 4082
rect 4558 4014 4698 4048
rect 4558 3980 4611 4014
rect 4645 3980 4698 4014
rect 4558 3946 4698 3980
rect 4558 3912 4611 3946
rect 4645 3912 4698 3946
rect 4558 3878 4698 3912
rect 4558 3844 4611 3878
rect 4645 3844 4698 3878
rect 4558 3810 4698 3844
rect 4558 3776 4611 3810
rect 4645 3776 4698 3810
rect 4558 3742 4698 3776
rect 4558 3708 4611 3742
rect 4645 3708 4698 3742
rect 4558 3674 4698 3708
rect 4558 3640 4611 3674
rect 4645 3640 4698 3674
rect 4558 3606 4698 3640
rect 4558 3572 4611 3606
rect 4645 3572 4698 3606
rect 4558 3538 4698 3572
rect 4558 3504 4611 3538
rect 4645 3504 4698 3538
rect 4558 3470 4698 3504
rect 4558 3436 4611 3470
rect 4645 3436 4698 3470
rect 4558 3402 4698 3436
rect 4558 3368 4611 3402
rect 4645 3368 4698 3402
rect 4558 3334 4698 3368
rect 4558 3300 4611 3334
rect 4645 3300 4698 3334
rect 4558 3266 4698 3300
rect 4558 3232 4611 3266
rect 4645 3232 4698 3266
rect 4558 3198 4698 3232
rect 4558 3164 4611 3198
rect 4645 3164 4698 3198
rect 4558 3152 4698 3164
rect 5550 4082 5690 4152
rect 5550 4048 5603 4082
rect 5637 4048 5690 4082
rect 5550 4014 5690 4048
rect 5550 3980 5603 4014
rect 5637 3980 5690 4014
rect 5550 3946 5690 3980
rect 5550 3912 5603 3946
rect 5637 3912 5690 3946
rect 5550 3878 5690 3912
rect 5550 3844 5603 3878
rect 5637 3844 5690 3878
rect 5550 3810 5690 3844
rect 5550 3776 5603 3810
rect 5637 3776 5690 3810
rect 5550 3742 5690 3776
rect 5550 3708 5603 3742
rect 5637 3708 5690 3742
rect 5550 3674 5690 3708
rect 5550 3640 5603 3674
rect 5637 3640 5690 3674
rect 5550 3606 5690 3640
rect 5550 3572 5603 3606
rect 5637 3572 5690 3606
rect 5550 3538 5690 3572
rect 5550 3504 5603 3538
rect 5637 3504 5690 3538
rect 5550 3470 5690 3504
rect 5550 3436 5603 3470
rect 5637 3436 5690 3470
rect 5550 3402 5690 3436
rect 5550 3368 5603 3402
rect 5637 3368 5690 3402
rect 5550 3334 5690 3368
rect 5550 3300 5603 3334
rect 5637 3300 5690 3334
rect 5550 3266 5690 3300
rect 5550 3232 5603 3266
rect 5637 3232 5690 3266
rect 5550 3198 5690 3232
rect 5550 3164 5603 3198
rect 5637 3164 5690 3198
rect 5550 3152 5690 3164
rect 6542 4082 6682 4152
rect 6542 4048 6595 4082
rect 6629 4048 6682 4082
rect 6542 4014 6682 4048
rect 6542 3980 6595 4014
rect 6629 3980 6682 4014
rect 6542 3946 6682 3980
rect 6542 3912 6595 3946
rect 6629 3912 6682 3946
rect 6542 3878 6682 3912
rect 6542 3844 6595 3878
rect 6629 3844 6682 3878
rect 6542 3810 6682 3844
rect 6542 3776 6595 3810
rect 6629 3776 6682 3810
rect 6542 3742 6682 3776
rect 6542 3708 6595 3742
rect 6629 3708 6682 3742
rect 6542 3674 6682 3708
rect 6542 3640 6595 3674
rect 6629 3640 6682 3674
rect 6542 3606 6682 3640
rect 6542 3572 6595 3606
rect 6629 3572 6682 3606
rect 6542 3538 6682 3572
rect 6542 3504 6595 3538
rect 6629 3504 6682 3538
rect 6542 3470 6682 3504
rect 6542 3436 6595 3470
rect 6629 3436 6682 3470
rect 6542 3402 6682 3436
rect 6542 3368 6595 3402
rect 6629 3368 6682 3402
rect 6542 3334 6682 3368
rect 6542 3300 6595 3334
rect 6629 3300 6682 3334
rect 6542 3266 6682 3300
rect 6542 3232 6595 3266
rect 6629 3232 6682 3266
rect 6542 3198 6682 3232
rect 6542 3164 6595 3198
rect 6629 3164 6682 3198
rect 6542 3152 6682 3164
rect 7534 4082 7674 4152
rect 7534 4048 7587 4082
rect 7621 4048 7674 4082
rect 7534 4014 7674 4048
rect 7534 3980 7587 4014
rect 7621 3980 7674 4014
rect 7534 3946 7674 3980
rect 7534 3912 7587 3946
rect 7621 3912 7674 3946
rect 7534 3878 7674 3912
rect 7534 3844 7587 3878
rect 7621 3844 7674 3878
rect 7534 3810 7674 3844
rect 7534 3776 7587 3810
rect 7621 3776 7674 3810
rect 7534 3742 7674 3776
rect 7534 3708 7587 3742
rect 7621 3708 7674 3742
rect 7534 3674 7674 3708
rect 7534 3640 7587 3674
rect 7621 3640 7674 3674
rect 7534 3606 7674 3640
rect 7534 3572 7587 3606
rect 7621 3572 7674 3606
rect 7534 3538 7674 3572
rect 7534 3504 7587 3538
rect 7621 3504 7674 3538
rect 7534 3470 7674 3504
rect 7534 3436 7587 3470
rect 7621 3436 7674 3470
rect 7534 3402 7674 3436
rect 7534 3368 7587 3402
rect 7621 3368 7674 3402
rect 7534 3334 7674 3368
rect 7534 3300 7587 3334
rect 7621 3300 7674 3334
rect 7534 3266 7674 3300
rect 7534 3232 7587 3266
rect 7621 3232 7674 3266
rect 7534 3198 7674 3232
rect 7534 3164 7587 3198
rect 7621 3164 7674 3198
rect 7534 3152 7674 3164
rect 8526 4082 8666 4152
rect 8526 4048 8579 4082
rect 8613 4048 8666 4082
rect 8526 4014 8666 4048
rect 8526 3980 8579 4014
rect 8613 3980 8666 4014
rect 8526 3946 8666 3980
rect 8526 3912 8579 3946
rect 8613 3912 8666 3946
rect 8526 3878 8666 3912
rect 8526 3844 8579 3878
rect 8613 3844 8666 3878
rect 8526 3810 8666 3844
rect 8526 3776 8579 3810
rect 8613 3776 8666 3810
rect 8526 3742 8666 3776
rect 8526 3708 8579 3742
rect 8613 3708 8666 3742
rect 8526 3674 8666 3708
rect 8526 3640 8579 3674
rect 8613 3640 8666 3674
rect 8526 3606 8666 3640
rect 8526 3572 8579 3606
rect 8613 3572 8666 3606
rect 8526 3538 8666 3572
rect 8526 3504 8579 3538
rect 8613 3504 8666 3538
rect 8526 3470 8666 3504
rect 8526 3436 8579 3470
rect 8613 3436 8666 3470
rect 8526 3402 8666 3436
rect 8526 3368 8579 3402
rect 8613 3368 8666 3402
rect 8526 3334 8666 3368
rect 8526 3300 8579 3334
rect 8613 3300 8666 3334
rect 8526 3266 8666 3300
rect 8526 3232 8579 3266
rect 8613 3232 8666 3266
rect 8526 3198 8666 3232
rect 8526 3164 8579 3198
rect 8613 3164 8666 3198
rect 8526 3152 8666 3164
rect 9518 4082 9658 4152
rect 9518 4048 9571 4082
rect 9605 4048 9658 4082
rect 9518 4014 9658 4048
rect 9518 3980 9571 4014
rect 9605 3980 9658 4014
rect 9518 3946 9658 3980
rect 9518 3912 9571 3946
rect 9605 3912 9658 3946
rect 9518 3878 9658 3912
rect 9518 3844 9571 3878
rect 9605 3844 9658 3878
rect 9518 3810 9658 3844
rect 9518 3776 9571 3810
rect 9605 3776 9658 3810
rect 9518 3742 9658 3776
rect 9518 3708 9571 3742
rect 9605 3708 9658 3742
rect 9518 3674 9658 3708
rect 9518 3640 9571 3674
rect 9605 3640 9658 3674
rect 9518 3606 9658 3640
rect 9518 3572 9571 3606
rect 9605 3572 9658 3606
rect 9518 3538 9658 3572
rect 9518 3504 9571 3538
rect 9605 3504 9658 3538
rect 9518 3470 9658 3504
rect 9518 3436 9571 3470
rect 9605 3436 9658 3470
rect 9518 3402 9658 3436
rect 9518 3368 9571 3402
rect 9605 3368 9658 3402
rect 9518 3334 9658 3368
rect 9518 3300 9571 3334
rect 9605 3300 9658 3334
rect 9518 3266 9658 3300
rect 9518 3232 9571 3266
rect 9605 3232 9658 3266
rect 9518 3198 9658 3232
rect 9518 3164 9571 3198
rect 9605 3164 9658 3198
rect 9518 3152 9658 3164
rect 10510 4082 10650 4152
rect 10510 4048 10563 4082
rect 10597 4048 10650 4082
rect 10510 4014 10650 4048
rect 10510 3980 10563 4014
rect 10597 3980 10650 4014
rect 10510 3946 10650 3980
rect 10510 3912 10563 3946
rect 10597 3912 10650 3946
rect 10510 3878 10650 3912
rect 10510 3844 10563 3878
rect 10597 3844 10650 3878
rect 10510 3810 10650 3844
rect 10510 3776 10563 3810
rect 10597 3776 10650 3810
rect 10510 3742 10650 3776
rect 10510 3708 10563 3742
rect 10597 3708 10650 3742
rect 10510 3674 10650 3708
rect 10510 3640 10563 3674
rect 10597 3640 10650 3674
rect 10510 3606 10650 3640
rect 10510 3572 10563 3606
rect 10597 3572 10650 3606
rect 10510 3538 10650 3572
rect 10510 3504 10563 3538
rect 10597 3504 10650 3538
rect 10510 3470 10650 3504
rect 10510 3436 10563 3470
rect 10597 3436 10650 3470
rect 10510 3402 10650 3436
rect 10510 3368 10563 3402
rect 10597 3368 10650 3402
rect 10510 3334 10650 3368
rect 10510 3300 10563 3334
rect 10597 3300 10650 3334
rect 10510 3266 10650 3300
rect 10510 3232 10563 3266
rect 10597 3232 10650 3266
rect 10510 3198 10650 3232
rect 10510 3164 10563 3198
rect 10597 3164 10650 3198
rect 10510 3152 10650 3164
rect 11502 4082 11642 4152
rect 11502 4048 11555 4082
rect 11589 4048 11642 4082
rect 11502 4014 11642 4048
rect 11502 3980 11555 4014
rect 11589 3980 11642 4014
rect 11502 3946 11642 3980
rect 11502 3912 11555 3946
rect 11589 3912 11642 3946
rect 11502 3878 11642 3912
rect 11502 3844 11555 3878
rect 11589 3844 11642 3878
rect 11502 3810 11642 3844
rect 11502 3776 11555 3810
rect 11589 3776 11642 3810
rect 11502 3742 11642 3776
rect 11502 3708 11555 3742
rect 11589 3708 11642 3742
rect 11502 3674 11642 3708
rect 11502 3640 11555 3674
rect 11589 3640 11642 3674
rect 11502 3606 11642 3640
rect 11502 3572 11555 3606
rect 11589 3572 11642 3606
rect 11502 3538 11642 3572
rect 11502 3504 11555 3538
rect 11589 3504 11642 3538
rect 11502 3470 11642 3504
rect 11502 3436 11555 3470
rect 11589 3436 11642 3470
rect 11502 3402 11642 3436
rect 11502 3368 11555 3402
rect 11589 3368 11642 3402
rect 11502 3334 11642 3368
rect 11502 3300 11555 3334
rect 11589 3300 11642 3334
rect 11502 3266 11642 3300
rect 11502 3232 11555 3266
rect 11589 3232 11642 3266
rect 11502 3198 11642 3232
rect 11502 3164 11555 3198
rect 11589 3164 11642 3198
rect 11502 3152 11642 3164
rect 12494 4082 12634 4152
rect 12494 4048 12547 4082
rect 12581 4048 12634 4082
rect 12494 4014 12634 4048
rect 12494 3980 12547 4014
rect 12581 3980 12634 4014
rect 12494 3946 12634 3980
rect 12494 3912 12547 3946
rect 12581 3912 12634 3946
rect 12494 3878 12634 3912
rect 12494 3844 12547 3878
rect 12581 3844 12634 3878
rect 12494 3810 12634 3844
rect 12494 3776 12547 3810
rect 12581 3776 12634 3810
rect 12494 3742 12634 3776
rect 12494 3708 12547 3742
rect 12581 3708 12634 3742
rect 12494 3674 12634 3708
rect 12494 3640 12547 3674
rect 12581 3640 12634 3674
rect 12494 3606 12634 3640
rect 12494 3572 12547 3606
rect 12581 3572 12634 3606
rect 12494 3538 12634 3572
rect 12494 3504 12547 3538
rect 12581 3504 12634 3538
rect 12494 3470 12634 3504
rect 12494 3436 12547 3470
rect 12581 3436 12634 3470
rect 12494 3402 12634 3436
rect 12494 3368 12547 3402
rect 12581 3368 12634 3402
rect 12494 3334 12634 3368
rect 12494 3300 12547 3334
rect 12581 3300 12634 3334
rect 12494 3266 12634 3300
rect 12494 3232 12547 3266
rect 12581 3232 12634 3266
rect 12494 3198 12634 3232
rect 12494 3164 12547 3198
rect 12581 3164 12634 3198
rect 12494 3152 12634 3164
rect 13486 4082 13626 4152
rect 13486 4048 13539 4082
rect 13573 4048 13626 4082
rect 13486 4014 13626 4048
rect 13486 3980 13539 4014
rect 13573 3980 13626 4014
rect 13486 3946 13626 3980
rect 13486 3912 13539 3946
rect 13573 3912 13626 3946
rect 13486 3878 13626 3912
rect 13486 3844 13539 3878
rect 13573 3844 13626 3878
rect 13486 3810 13626 3844
rect 13486 3776 13539 3810
rect 13573 3776 13626 3810
rect 13486 3742 13626 3776
rect 13486 3708 13539 3742
rect 13573 3708 13626 3742
rect 13486 3674 13626 3708
rect 13486 3640 13539 3674
rect 13573 3640 13626 3674
rect 13486 3606 13626 3640
rect 13486 3572 13539 3606
rect 13573 3572 13626 3606
rect 13486 3538 13626 3572
rect 13486 3504 13539 3538
rect 13573 3504 13626 3538
rect 13486 3470 13626 3504
rect 13486 3436 13539 3470
rect 13573 3436 13626 3470
rect 13486 3402 13626 3436
rect 13486 3368 13539 3402
rect 13573 3368 13626 3402
rect 13486 3334 13626 3368
rect 13486 3300 13539 3334
rect 13573 3300 13626 3334
rect 13486 3266 13626 3300
rect 13486 3232 13539 3266
rect 13573 3232 13626 3266
rect 13486 3198 13626 3232
rect 13486 3164 13539 3198
rect 13573 3164 13626 3198
rect 13486 3152 13626 3164
rect 14427 3992 14468 4152
rect 14427 3957 14536 3992
rect 14427 3923 14468 3957
rect 14502 3924 14536 3957
rect 14502 3923 14604 3924
rect 14427 3905 14604 3923
rect 14638 3905 14653 4551
rect 14427 3889 14653 3905
rect 14427 3888 14536 3889
rect 14427 3854 14468 3888
rect 14502 3855 14536 3888
rect 14570 3871 14653 3889
rect 14570 3855 14604 3871
rect 14502 3854 14604 3855
rect 14427 3837 14604 3854
rect 14638 3837 14653 3871
rect 14427 3820 14653 3837
rect 14427 3819 14536 3820
rect 14427 3785 14468 3819
rect 14502 3786 14536 3819
rect 14570 3803 14653 3820
rect 14570 3786 14604 3803
rect 14502 3785 14604 3786
rect 14427 3769 14604 3785
rect 14638 3769 14653 3803
rect 14427 3751 14653 3769
rect 14427 3750 14536 3751
rect 14427 3716 14468 3750
rect 14502 3717 14536 3750
rect 14570 3735 14653 3751
rect 14570 3717 14604 3735
rect 14502 3716 14604 3717
rect 14427 3701 14604 3716
rect 14638 3701 14653 3735
rect 14427 3682 14653 3701
rect 14427 3681 14536 3682
rect 14427 3647 14468 3681
rect 14502 3648 14536 3681
rect 14570 3667 14653 3682
rect 14570 3648 14604 3667
rect 14502 3647 14604 3648
rect 14427 3633 14604 3647
rect 14638 3633 14653 3667
rect 14427 3613 14653 3633
rect 14427 3612 14536 3613
rect 14427 3578 14468 3612
rect 14502 3579 14536 3612
rect 14570 3599 14653 3613
rect 14570 3579 14604 3599
rect 14502 3578 14604 3579
rect 14427 3565 14604 3578
rect 14638 3565 14653 3599
rect 14427 3544 14653 3565
rect 14427 3543 14536 3544
rect 14427 3509 14468 3543
rect 14502 3510 14536 3543
rect 14570 3531 14653 3544
rect 14570 3510 14604 3531
rect 14502 3509 14604 3510
rect 14427 3497 14604 3509
rect 14638 3497 14653 3531
rect 14427 3475 14653 3497
rect 14427 3474 14536 3475
rect 14427 3440 14468 3474
rect 14502 3441 14536 3474
rect 14570 3463 14653 3475
rect 14570 3441 14604 3463
rect 14502 3440 14604 3441
rect 14427 3429 14604 3440
rect 14638 3429 14653 3463
rect 14427 3406 14653 3429
rect 14427 3405 14536 3406
rect 14427 3371 14468 3405
rect 14502 3372 14536 3405
rect 14570 3395 14653 3406
rect 14570 3372 14604 3395
rect 14502 3371 14604 3372
rect 14427 3361 14604 3371
rect 14638 3361 14653 3395
rect 14427 3337 14653 3361
rect 14427 3336 14536 3337
rect 14427 3302 14468 3336
rect 14502 3303 14536 3336
rect 14570 3327 14653 3337
rect 14570 3303 14604 3327
rect 14502 3302 14604 3303
rect 14427 3293 14604 3302
rect 14638 3293 14653 3327
rect 14427 3268 14653 3293
rect 14427 3267 14536 3268
rect 14427 3233 14468 3267
rect 14502 3234 14536 3267
rect 14570 3259 14653 3268
rect 14570 3234 14604 3259
rect 14502 3233 14604 3234
rect 14427 3225 14604 3233
rect 14638 3225 14653 3259
rect 14427 3199 14653 3225
rect 14427 3198 14536 3199
rect 14427 3164 14468 3198
rect 14502 3165 14536 3198
rect 14570 3191 14653 3199
rect 14570 3165 14604 3191
rect 14502 3164 14604 3165
rect 14427 3157 14604 3164
rect 14638 3157 14653 3191
rect 14427 3152 14653 3157
rect 482 3128 682 3152
rect 482 3094 497 3128
rect 531 3094 565 3128
rect 599 3094 633 3128
rect 667 3094 682 3128
rect 482 3059 682 3094
rect 482 3025 497 3059
rect 531 3025 565 3059
rect 599 3025 633 3059
rect 667 3025 682 3059
rect 482 2990 682 3025
rect 482 2956 497 2990
rect 531 2956 565 2990
rect 599 2956 633 2990
rect 667 2956 682 2990
rect 482 2921 682 2956
rect 482 2887 497 2921
rect 531 2887 565 2921
rect 599 2887 633 2921
rect 667 2887 682 2921
rect 482 2852 682 2887
rect 482 2818 497 2852
rect 531 2818 565 2852
rect 599 2818 633 2852
rect 667 2818 682 2852
rect 482 2783 682 2818
rect 482 2749 497 2783
rect 531 2749 565 2783
rect 599 2749 633 2783
rect 667 2749 682 2783
rect 482 2714 682 2749
rect 482 2680 497 2714
rect 531 2680 565 2714
rect 599 2680 633 2714
rect 667 2680 682 2714
rect 482 2645 682 2680
rect 482 2611 497 2645
rect 531 2611 565 2645
rect 599 2611 633 2645
rect 667 2611 682 2645
rect 482 2576 682 2611
rect 482 2542 497 2576
rect 531 2542 565 2576
rect 599 2542 633 2576
rect 667 2552 682 2576
rect 1541 3044 1763 3078
rect 1541 3010 1601 3044
rect 1635 3010 1669 3044
rect 1703 3010 1763 3044
rect 1541 2974 1763 3010
rect 1541 2940 1601 2974
rect 1635 2940 1669 2974
rect 1703 2940 1763 2974
rect 1541 2904 1763 2940
rect 1541 2870 1601 2904
rect 1635 2870 1669 2904
rect 1703 2870 1763 2904
rect 1541 2834 1763 2870
rect 1541 2800 1601 2834
rect 1635 2800 1669 2834
rect 1703 2800 1763 2834
rect 1541 2764 1763 2800
rect 1541 2730 1601 2764
rect 1635 2730 1669 2764
rect 1703 2730 1763 2764
rect 1541 2694 1763 2730
rect 1541 2660 1601 2694
rect 1635 2660 1669 2694
rect 1703 2660 1763 2694
rect 1541 2626 1763 2660
rect 2533 3044 2755 3078
rect 2533 3010 2593 3044
rect 2627 3010 2661 3044
rect 2695 3010 2755 3044
rect 2533 2974 2755 3010
rect 2533 2940 2593 2974
rect 2627 2940 2661 2974
rect 2695 2940 2755 2974
rect 2533 2904 2755 2940
rect 2533 2870 2593 2904
rect 2627 2870 2661 2904
rect 2695 2870 2755 2904
rect 2533 2834 2755 2870
rect 2533 2800 2593 2834
rect 2627 2800 2661 2834
rect 2695 2800 2755 2834
rect 2533 2764 2755 2800
rect 2533 2730 2593 2764
rect 2627 2730 2661 2764
rect 2695 2730 2755 2764
rect 2533 2694 2755 2730
rect 2533 2660 2593 2694
rect 2627 2660 2661 2694
rect 2695 2660 2755 2694
rect 2533 2626 2755 2660
rect 3525 3044 3747 3078
rect 3525 3010 3585 3044
rect 3619 3010 3653 3044
rect 3687 3010 3747 3044
rect 3525 2974 3747 3010
rect 3525 2940 3585 2974
rect 3619 2940 3653 2974
rect 3687 2940 3747 2974
rect 3525 2904 3747 2940
rect 3525 2870 3585 2904
rect 3619 2870 3653 2904
rect 3687 2870 3747 2904
rect 3525 2834 3747 2870
rect 3525 2800 3585 2834
rect 3619 2800 3653 2834
rect 3687 2800 3747 2834
rect 3525 2764 3747 2800
rect 3525 2730 3585 2764
rect 3619 2730 3653 2764
rect 3687 2730 3747 2764
rect 3525 2694 3747 2730
rect 3525 2660 3585 2694
rect 3619 2660 3653 2694
rect 3687 2660 3747 2694
rect 3525 2626 3747 2660
rect 4517 3044 4739 3078
rect 4517 3010 4577 3044
rect 4611 3010 4645 3044
rect 4679 3010 4739 3044
rect 4517 2974 4739 3010
rect 4517 2940 4577 2974
rect 4611 2940 4645 2974
rect 4679 2940 4739 2974
rect 4517 2904 4739 2940
rect 4517 2870 4577 2904
rect 4611 2870 4645 2904
rect 4679 2870 4739 2904
rect 4517 2834 4739 2870
rect 4517 2800 4577 2834
rect 4611 2800 4645 2834
rect 4679 2800 4739 2834
rect 4517 2764 4739 2800
rect 4517 2730 4577 2764
rect 4611 2730 4645 2764
rect 4679 2730 4739 2764
rect 4517 2694 4739 2730
rect 4517 2660 4577 2694
rect 4611 2660 4645 2694
rect 4679 2660 4739 2694
rect 4517 2626 4739 2660
rect 5509 3044 5731 3078
rect 5509 3010 5569 3044
rect 5603 3010 5637 3044
rect 5671 3010 5731 3044
rect 5509 2974 5731 3010
rect 5509 2940 5569 2974
rect 5603 2940 5637 2974
rect 5671 2940 5731 2974
rect 5509 2904 5731 2940
rect 5509 2870 5569 2904
rect 5603 2870 5637 2904
rect 5671 2870 5731 2904
rect 5509 2834 5731 2870
rect 5509 2800 5569 2834
rect 5603 2800 5637 2834
rect 5671 2800 5731 2834
rect 5509 2764 5731 2800
rect 5509 2730 5569 2764
rect 5603 2730 5637 2764
rect 5671 2730 5731 2764
rect 5509 2694 5731 2730
rect 5509 2660 5569 2694
rect 5603 2660 5637 2694
rect 5671 2660 5731 2694
rect 5509 2626 5731 2660
rect 6501 3044 6723 3078
rect 6501 3010 6561 3044
rect 6595 3010 6629 3044
rect 6663 3010 6723 3044
rect 6501 2974 6723 3010
rect 6501 2940 6561 2974
rect 6595 2940 6629 2974
rect 6663 2940 6723 2974
rect 6501 2904 6723 2940
rect 6501 2870 6561 2904
rect 6595 2870 6629 2904
rect 6663 2870 6723 2904
rect 6501 2834 6723 2870
rect 6501 2800 6561 2834
rect 6595 2800 6629 2834
rect 6663 2800 6723 2834
rect 6501 2764 6723 2800
rect 6501 2730 6561 2764
rect 6595 2730 6629 2764
rect 6663 2730 6723 2764
rect 6501 2694 6723 2730
rect 6501 2660 6561 2694
rect 6595 2660 6629 2694
rect 6663 2660 6723 2694
rect 6501 2626 6723 2660
rect 7493 3044 7715 3078
rect 7493 3010 7553 3044
rect 7587 3010 7621 3044
rect 7655 3010 7715 3044
rect 7493 2974 7715 3010
rect 7493 2940 7553 2974
rect 7587 2940 7621 2974
rect 7655 2940 7715 2974
rect 7493 2904 7715 2940
rect 7493 2870 7553 2904
rect 7587 2870 7621 2904
rect 7655 2870 7715 2904
rect 7493 2834 7715 2870
rect 7493 2800 7553 2834
rect 7587 2800 7621 2834
rect 7655 2800 7715 2834
rect 7493 2764 7715 2800
rect 7493 2730 7553 2764
rect 7587 2730 7621 2764
rect 7655 2730 7715 2764
rect 7493 2694 7715 2730
rect 7493 2660 7553 2694
rect 7587 2660 7621 2694
rect 7655 2660 7715 2694
rect 7493 2626 7715 2660
rect 8485 3044 8707 3078
rect 8485 3010 8545 3044
rect 8579 3010 8613 3044
rect 8647 3010 8707 3044
rect 8485 2974 8707 3010
rect 8485 2940 8545 2974
rect 8579 2940 8613 2974
rect 8647 2940 8707 2974
rect 8485 2904 8707 2940
rect 8485 2870 8545 2904
rect 8579 2870 8613 2904
rect 8647 2870 8707 2904
rect 8485 2834 8707 2870
rect 8485 2800 8545 2834
rect 8579 2800 8613 2834
rect 8647 2800 8707 2834
rect 8485 2764 8707 2800
rect 8485 2730 8545 2764
rect 8579 2730 8613 2764
rect 8647 2730 8707 2764
rect 8485 2694 8707 2730
rect 8485 2660 8545 2694
rect 8579 2660 8613 2694
rect 8647 2660 8707 2694
rect 8485 2626 8707 2660
rect 9477 3044 9699 3078
rect 9477 3010 9537 3044
rect 9571 3010 9605 3044
rect 9639 3010 9699 3044
rect 9477 2974 9699 3010
rect 9477 2940 9537 2974
rect 9571 2940 9605 2974
rect 9639 2940 9699 2974
rect 9477 2904 9699 2940
rect 9477 2870 9537 2904
rect 9571 2870 9605 2904
rect 9639 2870 9699 2904
rect 9477 2834 9699 2870
rect 9477 2800 9537 2834
rect 9571 2800 9605 2834
rect 9639 2800 9699 2834
rect 9477 2764 9699 2800
rect 9477 2730 9537 2764
rect 9571 2730 9605 2764
rect 9639 2730 9699 2764
rect 9477 2694 9699 2730
rect 9477 2660 9537 2694
rect 9571 2660 9605 2694
rect 9639 2660 9699 2694
rect 9477 2626 9699 2660
rect 10469 3044 10691 3078
rect 10469 3010 10529 3044
rect 10563 3010 10597 3044
rect 10631 3010 10691 3044
rect 10469 2974 10691 3010
rect 10469 2940 10529 2974
rect 10563 2940 10597 2974
rect 10631 2940 10691 2974
rect 10469 2904 10691 2940
rect 10469 2870 10529 2904
rect 10563 2870 10597 2904
rect 10631 2870 10691 2904
rect 10469 2834 10691 2870
rect 10469 2800 10529 2834
rect 10563 2800 10597 2834
rect 10631 2800 10691 2834
rect 10469 2764 10691 2800
rect 10469 2730 10529 2764
rect 10563 2730 10597 2764
rect 10631 2730 10691 2764
rect 10469 2694 10691 2730
rect 10469 2660 10529 2694
rect 10563 2660 10597 2694
rect 10631 2660 10691 2694
rect 10469 2626 10691 2660
rect 11461 3044 11683 3078
rect 11461 3010 11521 3044
rect 11555 3010 11589 3044
rect 11623 3010 11683 3044
rect 11461 2974 11683 3010
rect 11461 2940 11521 2974
rect 11555 2940 11589 2974
rect 11623 2940 11683 2974
rect 11461 2904 11683 2940
rect 11461 2870 11521 2904
rect 11555 2870 11589 2904
rect 11623 2870 11683 2904
rect 11461 2834 11683 2870
rect 11461 2800 11521 2834
rect 11555 2800 11589 2834
rect 11623 2800 11683 2834
rect 11461 2764 11683 2800
rect 11461 2730 11521 2764
rect 11555 2730 11589 2764
rect 11623 2730 11683 2764
rect 11461 2694 11683 2730
rect 11461 2660 11521 2694
rect 11555 2660 11589 2694
rect 11623 2660 11683 2694
rect 11461 2626 11683 2660
rect 12453 3044 12675 3078
rect 12453 3010 12513 3044
rect 12547 3010 12581 3044
rect 12615 3010 12675 3044
rect 12453 2974 12675 3010
rect 12453 2940 12513 2974
rect 12547 2940 12581 2974
rect 12615 2940 12675 2974
rect 12453 2904 12675 2940
rect 12453 2870 12513 2904
rect 12547 2870 12581 2904
rect 12615 2870 12675 2904
rect 12453 2834 12675 2870
rect 12453 2800 12513 2834
rect 12547 2800 12581 2834
rect 12615 2800 12675 2834
rect 12453 2764 12675 2800
rect 12453 2730 12513 2764
rect 12547 2730 12581 2764
rect 12615 2730 12675 2764
rect 12453 2694 12675 2730
rect 12453 2660 12513 2694
rect 12547 2660 12581 2694
rect 12615 2660 12675 2694
rect 12453 2626 12675 2660
rect 13445 3044 13667 3078
rect 13445 3010 13505 3044
rect 13539 3010 13573 3044
rect 13607 3010 13667 3044
rect 13445 2974 13667 3010
rect 13445 2940 13505 2974
rect 13539 2940 13573 2974
rect 13607 2940 13667 2974
rect 13445 2904 13667 2940
rect 13445 2870 13505 2904
rect 13539 2870 13573 2904
rect 13607 2870 13667 2904
rect 13445 2834 13667 2870
rect 13445 2800 13505 2834
rect 13539 2800 13573 2834
rect 13607 2800 13667 2834
rect 13445 2764 13667 2800
rect 13445 2730 13505 2764
rect 13539 2730 13573 2764
rect 13607 2730 13667 2764
rect 13445 2694 13667 2730
rect 13445 2660 13505 2694
rect 13539 2660 13573 2694
rect 13607 2660 13667 2694
rect 13445 2626 13667 2660
rect 14453 3130 14653 3152
rect 14453 3129 14536 3130
rect 14453 3095 14468 3129
rect 14502 3096 14536 3129
rect 14570 3123 14653 3130
rect 14570 3096 14604 3123
rect 14502 3095 14604 3096
rect 14453 3089 14604 3095
rect 14638 3089 14653 3123
rect 14453 3061 14653 3089
rect 14453 3060 14536 3061
rect 14453 3026 14468 3060
rect 14502 3027 14536 3060
rect 14570 3055 14653 3061
rect 14570 3027 14604 3055
rect 14502 3026 14604 3027
rect 14453 3021 14604 3026
rect 14638 3021 14653 3055
rect 14453 2992 14653 3021
rect 14453 2991 14536 2992
rect 14453 2957 14468 2991
rect 14502 2958 14536 2991
rect 14570 2987 14653 2992
rect 14570 2958 14604 2987
rect 14502 2957 14604 2958
rect 14453 2953 14604 2957
rect 14638 2953 14653 2987
rect 14453 2923 14653 2953
rect 14453 2922 14536 2923
rect 14453 2888 14468 2922
rect 14502 2889 14536 2922
rect 14570 2919 14653 2923
rect 14570 2889 14604 2919
rect 14502 2888 14604 2889
rect 14453 2885 14604 2888
rect 14638 2885 14653 2919
rect 14453 2854 14653 2885
rect 14453 2853 14536 2854
rect 14453 2819 14468 2853
rect 14502 2820 14536 2853
rect 14570 2851 14653 2854
rect 14570 2820 14604 2851
rect 14502 2819 14604 2820
rect 14453 2817 14604 2819
rect 14638 2817 14653 2851
rect 14453 2785 14653 2817
rect 14453 2784 14536 2785
rect 14453 2750 14468 2784
rect 14502 2751 14536 2784
rect 14570 2783 14653 2785
rect 14570 2751 14604 2783
rect 14502 2750 14604 2751
rect 14453 2749 14604 2750
rect 14638 2749 14653 2783
rect 14453 2716 14653 2749
rect 14453 2715 14536 2716
rect 14453 2681 14468 2715
rect 14502 2682 14536 2715
rect 14570 2715 14653 2716
rect 14570 2682 14604 2715
rect 14502 2681 14604 2682
rect 14638 2681 14653 2715
rect 14453 2647 14653 2681
rect 14453 2646 14536 2647
rect 14453 2612 14468 2646
rect 14502 2613 14536 2646
rect 14570 2613 14604 2647
rect 14638 2613 14653 2647
rect 14502 2612 14653 2613
rect 14453 2579 14653 2612
rect 14453 2578 14604 2579
rect 14453 2577 14536 2578
rect 14453 2552 14468 2577
rect 667 2542 708 2552
rect 482 2507 708 2542
rect 482 2473 497 2507
rect 531 2473 565 2507
rect 599 2473 633 2507
rect 667 2473 708 2507
rect 482 2438 708 2473
rect 482 2404 497 2438
rect 531 2404 565 2438
rect 599 2404 633 2438
rect 667 2404 708 2438
rect 482 2369 708 2404
rect 482 2335 497 2369
rect 531 2335 565 2369
rect 599 2335 633 2369
rect 667 2335 708 2369
rect 482 2300 708 2335
rect 482 2266 497 2300
rect 531 2266 565 2300
rect 599 2266 633 2300
rect 667 2266 708 2300
rect 482 2231 708 2266
rect 482 2197 497 2231
rect 531 2197 565 2231
rect 599 2197 633 2231
rect 667 2197 708 2231
rect 482 2163 708 2197
rect 482 2129 497 2163
rect 531 2162 708 2163
rect 531 2129 565 2162
rect 482 2128 565 2129
rect 599 2128 633 2162
rect 667 2128 708 2162
rect 482 2095 708 2128
rect 482 2061 497 2095
rect 531 2093 708 2095
rect 531 2061 565 2093
rect 482 2059 565 2061
rect 599 2059 633 2093
rect 667 2059 708 2093
rect 482 2027 708 2059
rect 482 1993 497 2027
rect 531 2024 708 2027
rect 531 1993 565 2024
rect 482 1990 565 1993
rect 599 1990 633 2024
rect 667 1990 708 2024
rect 482 1959 708 1990
rect 482 1925 497 1959
rect 531 1955 708 1959
rect 531 1925 565 1955
rect 482 1921 565 1925
rect 599 1921 633 1955
rect 667 1921 708 1955
rect 482 1891 708 1921
rect 482 1857 497 1891
rect 531 1886 708 1891
rect 531 1857 565 1886
rect 482 1852 565 1857
rect 599 1852 633 1886
rect 667 1852 708 1886
rect 482 1823 708 1852
rect 482 1789 497 1823
rect 531 1817 708 1823
rect 531 1789 565 1817
rect 482 1783 565 1789
rect 599 1783 633 1817
rect 667 1783 708 1817
rect 482 1755 708 1783
rect 482 1721 497 1755
rect 531 1748 708 1755
rect 531 1721 565 1748
rect 482 1714 565 1721
rect 599 1714 633 1748
rect 667 1714 708 1748
rect 482 1687 708 1714
rect 482 1653 497 1687
rect 531 1679 708 1687
rect 531 1653 565 1679
rect 482 1645 565 1653
rect 599 1645 633 1679
rect 667 1645 708 1679
rect 482 1619 708 1645
rect 482 1585 497 1619
rect 531 1610 708 1619
rect 531 1585 565 1610
rect 482 1576 565 1585
rect 599 1576 633 1610
rect 667 1576 708 1610
rect 482 1552 708 1576
rect 1582 2540 1722 2552
rect 1582 2506 1635 2540
rect 1669 2506 1722 2540
rect 1582 2472 1722 2506
rect 1582 2438 1635 2472
rect 1669 2438 1722 2472
rect 1582 2404 1722 2438
rect 1582 2370 1635 2404
rect 1669 2370 1722 2404
rect 1582 2336 1722 2370
rect 1582 2302 1635 2336
rect 1669 2302 1722 2336
rect 1582 2268 1722 2302
rect 1582 2234 1635 2268
rect 1669 2234 1722 2268
rect 1582 2200 1722 2234
rect 1582 2166 1635 2200
rect 1669 2166 1722 2200
rect 1582 2132 1722 2166
rect 1582 2098 1635 2132
rect 1669 2098 1722 2132
rect 1582 2064 1722 2098
rect 1582 2030 1635 2064
rect 1669 2030 1722 2064
rect 1582 1996 1722 2030
rect 1582 1962 1635 1996
rect 1669 1962 1722 1996
rect 1582 1928 1722 1962
rect 1582 1894 1635 1928
rect 1669 1894 1722 1928
rect 1582 1860 1722 1894
rect 1582 1826 1635 1860
rect 1669 1826 1722 1860
rect 1582 1792 1722 1826
rect 1582 1758 1635 1792
rect 1669 1758 1722 1792
rect 1582 1724 1722 1758
rect 1582 1690 1635 1724
rect 1669 1690 1722 1724
rect 1582 1656 1722 1690
rect 1582 1622 1635 1656
rect 1669 1622 1722 1656
rect 1582 1552 1722 1622
rect 2574 2540 2714 2552
rect 2574 2506 2627 2540
rect 2661 2506 2714 2540
rect 2574 2472 2714 2506
rect 2574 2438 2627 2472
rect 2661 2438 2714 2472
rect 2574 2404 2714 2438
rect 2574 2370 2627 2404
rect 2661 2370 2714 2404
rect 2574 2336 2714 2370
rect 2574 2302 2627 2336
rect 2661 2302 2714 2336
rect 2574 2268 2714 2302
rect 2574 2234 2627 2268
rect 2661 2234 2714 2268
rect 2574 2200 2714 2234
rect 2574 2166 2627 2200
rect 2661 2166 2714 2200
rect 2574 2132 2714 2166
rect 2574 2098 2627 2132
rect 2661 2098 2714 2132
rect 2574 2064 2714 2098
rect 2574 2030 2627 2064
rect 2661 2030 2714 2064
rect 2574 1996 2714 2030
rect 2574 1962 2627 1996
rect 2661 1962 2714 1996
rect 2574 1928 2714 1962
rect 2574 1894 2627 1928
rect 2661 1894 2714 1928
rect 2574 1860 2714 1894
rect 2574 1826 2627 1860
rect 2661 1826 2714 1860
rect 2574 1792 2714 1826
rect 2574 1758 2627 1792
rect 2661 1758 2714 1792
rect 2574 1724 2714 1758
rect 2574 1690 2627 1724
rect 2661 1690 2714 1724
rect 2574 1656 2714 1690
rect 2574 1622 2627 1656
rect 2661 1622 2714 1656
rect 2574 1552 2714 1622
rect 3566 2540 3706 2552
rect 3566 2506 3619 2540
rect 3653 2506 3706 2540
rect 3566 2472 3706 2506
rect 3566 2438 3619 2472
rect 3653 2438 3706 2472
rect 3566 2404 3706 2438
rect 3566 2370 3619 2404
rect 3653 2370 3706 2404
rect 3566 2336 3706 2370
rect 3566 2302 3619 2336
rect 3653 2302 3706 2336
rect 3566 2268 3706 2302
rect 3566 2234 3619 2268
rect 3653 2234 3706 2268
rect 3566 2200 3706 2234
rect 3566 2166 3619 2200
rect 3653 2166 3706 2200
rect 3566 2132 3706 2166
rect 3566 2098 3619 2132
rect 3653 2098 3706 2132
rect 3566 2064 3706 2098
rect 3566 2030 3619 2064
rect 3653 2030 3706 2064
rect 3566 1996 3706 2030
rect 3566 1962 3619 1996
rect 3653 1962 3706 1996
rect 3566 1928 3706 1962
rect 3566 1894 3619 1928
rect 3653 1894 3706 1928
rect 3566 1860 3706 1894
rect 3566 1826 3619 1860
rect 3653 1826 3706 1860
rect 3566 1792 3706 1826
rect 3566 1758 3619 1792
rect 3653 1758 3706 1792
rect 3566 1724 3706 1758
rect 3566 1690 3619 1724
rect 3653 1690 3706 1724
rect 3566 1656 3706 1690
rect 3566 1622 3619 1656
rect 3653 1622 3706 1656
rect 3566 1552 3706 1622
rect 4558 2540 4698 2552
rect 4558 2506 4611 2540
rect 4645 2506 4698 2540
rect 4558 2472 4698 2506
rect 4558 2438 4611 2472
rect 4645 2438 4698 2472
rect 4558 2404 4698 2438
rect 4558 2370 4611 2404
rect 4645 2370 4698 2404
rect 4558 2336 4698 2370
rect 4558 2302 4611 2336
rect 4645 2302 4698 2336
rect 4558 2268 4698 2302
rect 4558 2234 4611 2268
rect 4645 2234 4698 2268
rect 4558 2200 4698 2234
rect 4558 2166 4611 2200
rect 4645 2166 4698 2200
rect 4558 2132 4698 2166
rect 4558 2098 4611 2132
rect 4645 2098 4698 2132
rect 4558 2064 4698 2098
rect 4558 2030 4611 2064
rect 4645 2030 4698 2064
rect 4558 1996 4698 2030
rect 4558 1962 4611 1996
rect 4645 1962 4698 1996
rect 4558 1928 4698 1962
rect 4558 1894 4611 1928
rect 4645 1894 4698 1928
rect 4558 1860 4698 1894
rect 4558 1826 4611 1860
rect 4645 1826 4698 1860
rect 4558 1792 4698 1826
rect 4558 1758 4611 1792
rect 4645 1758 4698 1792
rect 4558 1724 4698 1758
rect 4558 1690 4611 1724
rect 4645 1690 4698 1724
rect 4558 1656 4698 1690
rect 4558 1622 4611 1656
rect 4645 1622 4698 1656
rect 4558 1552 4698 1622
rect 5550 2540 5690 2552
rect 5550 2506 5603 2540
rect 5637 2506 5690 2540
rect 5550 2472 5690 2506
rect 5550 2438 5603 2472
rect 5637 2438 5690 2472
rect 5550 2404 5690 2438
rect 5550 2370 5603 2404
rect 5637 2370 5690 2404
rect 5550 2336 5690 2370
rect 5550 2302 5603 2336
rect 5637 2302 5690 2336
rect 5550 2268 5690 2302
rect 5550 2234 5603 2268
rect 5637 2234 5690 2268
rect 5550 2200 5690 2234
rect 5550 2166 5603 2200
rect 5637 2166 5690 2200
rect 5550 2132 5690 2166
rect 5550 2098 5603 2132
rect 5637 2098 5690 2132
rect 5550 2064 5690 2098
rect 5550 2030 5603 2064
rect 5637 2030 5690 2064
rect 5550 1996 5690 2030
rect 5550 1962 5603 1996
rect 5637 1962 5690 1996
rect 5550 1928 5690 1962
rect 5550 1894 5603 1928
rect 5637 1894 5690 1928
rect 5550 1860 5690 1894
rect 5550 1826 5603 1860
rect 5637 1826 5690 1860
rect 5550 1792 5690 1826
rect 5550 1758 5603 1792
rect 5637 1758 5690 1792
rect 5550 1724 5690 1758
rect 5550 1690 5603 1724
rect 5637 1690 5690 1724
rect 5550 1656 5690 1690
rect 5550 1622 5603 1656
rect 5637 1622 5690 1656
rect 5550 1552 5690 1622
rect 6542 2540 6682 2552
rect 6542 2506 6595 2540
rect 6629 2506 6682 2540
rect 6542 2472 6682 2506
rect 6542 2438 6595 2472
rect 6629 2438 6682 2472
rect 6542 2404 6682 2438
rect 6542 2370 6595 2404
rect 6629 2370 6682 2404
rect 6542 2336 6682 2370
rect 6542 2302 6595 2336
rect 6629 2302 6682 2336
rect 6542 2268 6682 2302
rect 6542 2234 6595 2268
rect 6629 2234 6682 2268
rect 6542 2200 6682 2234
rect 6542 2166 6595 2200
rect 6629 2166 6682 2200
rect 6542 2132 6682 2166
rect 6542 2098 6595 2132
rect 6629 2098 6682 2132
rect 6542 2064 6682 2098
rect 6542 2030 6595 2064
rect 6629 2030 6682 2064
rect 6542 1996 6682 2030
rect 6542 1962 6595 1996
rect 6629 1962 6682 1996
rect 6542 1928 6682 1962
rect 6542 1894 6595 1928
rect 6629 1894 6682 1928
rect 6542 1860 6682 1894
rect 6542 1826 6595 1860
rect 6629 1826 6682 1860
rect 6542 1792 6682 1826
rect 6542 1758 6595 1792
rect 6629 1758 6682 1792
rect 6542 1724 6682 1758
rect 6542 1690 6595 1724
rect 6629 1690 6682 1724
rect 6542 1656 6682 1690
rect 6542 1622 6595 1656
rect 6629 1622 6682 1656
rect 6542 1552 6682 1622
rect 7534 2540 7674 2552
rect 7534 2506 7587 2540
rect 7621 2506 7674 2540
rect 7534 2472 7674 2506
rect 7534 2438 7587 2472
rect 7621 2438 7674 2472
rect 7534 2404 7674 2438
rect 7534 2370 7587 2404
rect 7621 2370 7674 2404
rect 7534 2336 7674 2370
rect 7534 2302 7587 2336
rect 7621 2302 7674 2336
rect 7534 2268 7674 2302
rect 7534 2234 7587 2268
rect 7621 2234 7674 2268
rect 7534 2200 7674 2234
rect 7534 2166 7587 2200
rect 7621 2166 7674 2200
rect 7534 2132 7674 2166
rect 7534 2098 7587 2132
rect 7621 2098 7674 2132
rect 7534 2064 7674 2098
rect 7534 2030 7587 2064
rect 7621 2030 7674 2064
rect 7534 1996 7674 2030
rect 7534 1962 7587 1996
rect 7621 1962 7674 1996
rect 7534 1928 7674 1962
rect 7534 1894 7587 1928
rect 7621 1894 7674 1928
rect 7534 1860 7674 1894
rect 7534 1826 7587 1860
rect 7621 1826 7674 1860
rect 7534 1792 7674 1826
rect 7534 1758 7587 1792
rect 7621 1758 7674 1792
rect 7534 1724 7674 1758
rect 7534 1690 7587 1724
rect 7621 1690 7674 1724
rect 7534 1656 7674 1690
rect 7534 1622 7587 1656
rect 7621 1622 7674 1656
rect 7534 1552 7674 1622
rect 8526 2540 8666 2552
rect 8526 2506 8579 2540
rect 8613 2506 8666 2540
rect 8526 2472 8666 2506
rect 8526 2438 8579 2472
rect 8613 2438 8666 2472
rect 8526 2404 8666 2438
rect 8526 2370 8579 2404
rect 8613 2370 8666 2404
rect 8526 2336 8666 2370
rect 8526 2302 8579 2336
rect 8613 2302 8666 2336
rect 8526 2268 8666 2302
rect 8526 2234 8579 2268
rect 8613 2234 8666 2268
rect 8526 2200 8666 2234
rect 8526 2166 8579 2200
rect 8613 2166 8666 2200
rect 8526 2132 8666 2166
rect 8526 2098 8579 2132
rect 8613 2098 8666 2132
rect 8526 2064 8666 2098
rect 8526 2030 8579 2064
rect 8613 2030 8666 2064
rect 8526 1996 8666 2030
rect 8526 1962 8579 1996
rect 8613 1962 8666 1996
rect 8526 1928 8666 1962
rect 8526 1894 8579 1928
rect 8613 1894 8666 1928
rect 8526 1860 8666 1894
rect 8526 1826 8579 1860
rect 8613 1826 8666 1860
rect 8526 1792 8666 1826
rect 8526 1758 8579 1792
rect 8613 1758 8666 1792
rect 8526 1724 8666 1758
rect 8526 1690 8579 1724
rect 8613 1690 8666 1724
rect 8526 1656 8666 1690
rect 8526 1622 8579 1656
rect 8613 1622 8666 1656
rect 8526 1552 8666 1622
rect 9518 2540 9658 2552
rect 9518 2506 9571 2540
rect 9605 2506 9658 2540
rect 9518 2472 9658 2506
rect 9518 2438 9571 2472
rect 9605 2438 9658 2472
rect 9518 2404 9658 2438
rect 9518 2370 9571 2404
rect 9605 2370 9658 2404
rect 9518 2336 9658 2370
rect 9518 2302 9571 2336
rect 9605 2302 9658 2336
rect 9518 2268 9658 2302
rect 9518 2234 9571 2268
rect 9605 2234 9658 2268
rect 9518 2200 9658 2234
rect 9518 2166 9571 2200
rect 9605 2166 9658 2200
rect 9518 2132 9658 2166
rect 9518 2098 9571 2132
rect 9605 2098 9658 2132
rect 9518 2064 9658 2098
rect 9518 2030 9571 2064
rect 9605 2030 9658 2064
rect 9518 1996 9658 2030
rect 9518 1962 9571 1996
rect 9605 1962 9658 1996
rect 9518 1928 9658 1962
rect 9518 1894 9571 1928
rect 9605 1894 9658 1928
rect 9518 1860 9658 1894
rect 9518 1826 9571 1860
rect 9605 1826 9658 1860
rect 9518 1792 9658 1826
rect 9518 1758 9571 1792
rect 9605 1758 9658 1792
rect 9518 1724 9658 1758
rect 9518 1690 9571 1724
rect 9605 1690 9658 1724
rect 9518 1656 9658 1690
rect 9518 1622 9571 1656
rect 9605 1622 9658 1656
rect 9518 1552 9658 1622
rect 10510 2540 10650 2552
rect 10510 2506 10563 2540
rect 10597 2506 10650 2540
rect 10510 2472 10650 2506
rect 10510 2438 10563 2472
rect 10597 2438 10650 2472
rect 10510 2404 10650 2438
rect 10510 2370 10563 2404
rect 10597 2370 10650 2404
rect 10510 2336 10650 2370
rect 10510 2302 10563 2336
rect 10597 2302 10650 2336
rect 10510 2268 10650 2302
rect 10510 2234 10563 2268
rect 10597 2234 10650 2268
rect 10510 2200 10650 2234
rect 10510 2166 10563 2200
rect 10597 2166 10650 2200
rect 10510 2132 10650 2166
rect 10510 2098 10563 2132
rect 10597 2098 10650 2132
rect 10510 2064 10650 2098
rect 10510 2030 10563 2064
rect 10597 2030 10650 2064
rect 10510 1996 10650 2030
rect 10510 1962 10563 1996
rect 10597 1962 10650 1996
rect 10510 1928 10650 1962
rect 10510 1894 10563 1928
rect 10597 1894 10650 1928
rect 10510 1860 10650 1894
rect 10510 1826 10563 1860
rect 10597 1826 10650 1860
rect 10510 1792 10650 1826
rect 10510 1758 10563 1792
rect 10597 1758 10650 1792
rect 10510 1724 10650 1758
rect 10510 1690 10563 1724
rect 10597 1690 10650 1724
rect 10510 1656 10650 1690
rect 10510 1622 10563 1656
rect 10597 1622 10650 1656
rect 10510 1552 10650 1622
rect 11502 2540 11642 2552
rect 11502 2506 11555 2540
rect 11589 2506 11642 2540
rect 11502 2472 11642 2506
rect 11502 2438 11555 2472
rect 11589 2438 11642 2472
rect 11502 2404 11642 2438
rect 11502 2370 11555 2404
rect 11589 2370 11642 2404
rect 11502 2336 11642 2370
rect 11502 2302 11555 2336
rect 11589 2302 11642 2336
rect 11502 2268 11642 2302
rect 11502 2234 11555 2268
rect 11589 2234 11642 2268
rect 11502 2200 11642 2234
rect 11502 2166 11555 2200
rect 11589 2166 11642 2200
rect 11502 2132 11642 2166
rect 11502 2098 11555 2132
rect 11589 2098 11642 2132
rect 11502 2064 11642 2098
rect 11502 2030 11555 2064
rect 11589 2030 11642 2064
rect 11502 1996 11642 2030
rect 11502 1962 11555 1996
rect 11589 1962 11642 1996
rect 11502 1928 11642 1962
rect 11502 1894 11555 1928
rect 11589 1894 11642 1928
rect 11502 1860 11642 1894
rect 11502 1826 11555 1860
rect 11589 1826 11642 1860
rect 11502 1792 11642 1826
rect 11502 1758 11555 1792
rect 11589 1758 11642 1792
rect 11502 1724 11642 1758
rect 11502 1690 11555 1724
rect 11589 1690 11642 1724
rect 11502 1656 11642 1690
rect 11502 1622 11555 1656
rect 11589 1622 11642 1656
rect 11502 1552 11642 1622
rect 12494 2540 12634 2552
rect 12494 2506 12547 2540
rect 12581 2506 12634 2540
rect 12494 2472 12634 2506
rect 12494 2438 12547 2472
rect 12581 2438 12634 2472
rect 12494 2404 12634 2438
rect 12494 2370 12547 2404
rect 12581 2370 12634 2404
rect 12494 2336 12634 2370
rect 12494 2302 12547 2336
rect 12581 2302 12634 2336
rect 12494 2268 12634 2302
rect 12494 2234 12547 2268
rect 12581 2234 12634 2268
rect 12494 2200 12634 2234
rect 12494 2166 12547 2200
rect 12581 2166 12634 2200
rect 12494 2132 12634 2166
rect 12494 2098 12547 2132
rect 12581 2098 12634 2132
rect 12494 2064 12634 2098
rect 12494 2030 12547 2064
rect 12581 2030 12634 2064
rect 12494 1996 12634 2030
rect 12494 1962 12547 1996
rect 12581 1962 12634 1996
rect 12494 1928 12634 1962
rect 12494 1894 12547 1928
rect 12581 1894 12634 1928
rect 12494 1860 12634 1894
rect 12494 1826 12547 1860
rect 12581 1826 12634 1860
rect 12494 1792 12634 1826
rect 12494 1758 12547 1792
rect 12581 1758 12634 1792
rect 12494 1724 12634 1758
rect 12494 1690 12547 1724
rect 12581 1690 12634 1724
rect 12494 1656 12634 1690
rect 12494 1622 12547 1656
rect 12581 1622 12634 1656
rect 12494 1552 12634 1622
rect 13486 2540 13626 2552
rect 13486 2506 13539 2540
rect 13573 2506 13626 2540
rect 13486 2472 13626 2506
rect 13486 2438 13539 2472
rect 13573 2438 13626 2472
rect 13486 2404 13626 2438
rect 13486 2370 13539 2404
rect 13573 2370 13626 2404
rect 13486 2336 13626 2370
rect 13486 2302 13539 2336
rect 13573 2302 13626 2336
rect 13486 2268 13626 2302
rect 13486 2234 13539 2268
rect 13573 2234 13626 2268
rect 13486 2200 13626 2234
rect 13486 2166 13539 2200
rect 13573 2166 13626 2200
rect 13486 2132 13626 2166
rect 13486 2098 13539 2132
rect 13573 2098 13626 2132
rect 13486 2064 13626 2098
rect 13486 2030 13539 2064
rect 13573 2030 13626 2064
rect 13486 1996 13626 2030
rect 13486 1962 13539 1996
rect 13573 1962 13626 1996
rect 13486 1928 13626 1962
rect 13486 1894 13539 1928
rect 13573 1894 13626 1928
rect 13486 1860 13626 1894
rect 13486 1826 13539 1860
rect 13573 1826 13626 1860
rect 13486 1792 13626 1826
rect 13486 1758 13539 1792
rect 13573 1758 13626 1792
rect 13486 1724 13626 1758
rect 13486 1690 13539 1724
rect 13573 1690 13626 1724
rect 13486 1656 13626 1690
rect 13486 1622 13539 1656
rect 13573 1622 13626 1656
rect 13486 1552 13626 1622
rect 14427 2543 14468 2552
rect 14502 2544 14536 2577
rect 14570 2545 14604 2578
rect 14638 2545 14653 2579
rect 14570 2544 14653 2545
rect 14502 2543 14653 2544
rect 14427 2511 14653 2543
rect 14427 2509 14604 2511
rect 14427 2508 14536 2509
rect 14427 2474 14468 2508
rect 14502 2475 14536 2508
rect 14570 2477 14604 2509
rect 14638 2477 14653 2511
rect 14570 2475 14653 2477
rect 14502 2474 14653 2475
rect 14427 2443 14653 2474
rect 14427 2440 14604 2443
rect 14427 2439 14536 2440
rect 14427 2405 14468 2439
rect 14502 2406 14536 2439
rect 14570 2409 14604 2440
rect 14638 2409 14653 2443
rect 14570 2406 14653 2409
rect 14502 2405 14653 2406
rect 14427 2375 14653 2405
rect 14427 2371 14604 2375
rect 14427 2370 14536 2371
rect 14427 2336 14468 2370
rect 14502 2337 14536 2370
rect 14570 2341 14604 2371
rect 14638 2341 14653 2375
rect 14570 2337 14653 2341
rect 14502 2336 14653 2337
rect 14427 2307 14653 2336
rect 14427 2302 14604 2307
rect 14427 2301 14536 2302
rect 14427 2267 14468 2301
rect 14502 2268 14536 2301
rect 14570 2273 14604 2302
rect 14638 2273 14653 2307
rect 14570 2268 14653 2273
rect 14502 2267 14653 2268
rect 14427 2239 14653 2267
rect 14427 2233 14604 2239
rect 14427 2232 14536 2233
rect 14427 2198 14468 2232
rect 14502 2199 14536 2232
rect 14570 2205 14604 2233
rect 14638 2205 14653 2239
rect 14570 2199 14653 2205
rect 14502 2198 14653 2199
rect 14427 2171 14653 2198
rect 14427 2164 14604 2171
rect 14427 2163 14536 2164
rect 14427 2129 14468 2163
rect 14502 2130 14536 2163
rect 14570 2137 14604 2164
rect 14638 2137 14653 2171
rect 14570 2130 14653 2137
rect 14502 2129 14653 2130
rect 14427 2103 14653 2129
rect 14427 2095 14604 2103
rect 14427 2094 14536 2095
rect 14427 2060 14468 2094
rect 14502 2061 14536 2094
rect 14570 2069 14604 2095
rect 14638 2069 14653 2103
rect 14570 2061 14653 2069
rect 14502 2060 14653 2061
rect 14427 2035 14653 2060
rect 14427 2026 14604 2035
rect 14427 2025 14536 2026
rect 14427 1991 14468 2025
rect 14502 1992 14536 2025
rect 14570 2001 14604 2026
rect 14638 2001 14653 2035
rect 14570 1992 14653 2001
rect 14502 1991 14653 1992
rect 14427 1967 14653 1991
rect 14427 1957 14604 1967
rect 14427 1956 14536 1957
rect 14427 1922 14468 1956
rect 14502 1923 14536 1956
rect 14570 1933 14604 1957
rect 14638 1933 14653 1967
rect 14570 1923 14653 1933
rect 14502 1922 14653 1923
rect 14427 1899 14653 1922
rect 14427 1888 14604 1899
rect 14427 1887 14536 1888
rect 14427 1853 14468 1887
rect 14502 1854 14536 1887
rect 14570 1865 14604 1888
rect 14638 1865 14653 1899
rect 14570 1854 14653 1865
rect 14502 1853 14653 1854
rect 14427 1831 14653 1853
rect 14427 1819 14604 1831
rect 14427 1818 14536 1819
rect 14427 1784 14468 1818
rect 14502 1785 14536 1818
rect 14570 1797 14604 1819
rect 14638 1797 14653 1831
rect 14570 1785 14653 1797
rect 14502 1784 14653 1785
rect 14427 1763 14653 1784
rect 14427 1750 14604 1763
rect 14427 1749 14536 1750
rect 14427 1715 14468 1749
rect 14502 1716 14536 1749
rect 14570 1729 14604 1750
rect 14638 1729 14653 1763
rect 14570 1716 14653 1729
rect 14502 1715 14653 1716
rect 14427 1695 14653 1715
rect 14427 1681 14604 1695
rect 14427 1680 14536 1681
rect 14427 1646 14468 1680
rect 14502 1647 14536 1680
rect 14570 1661 14604 1681
rect 14638 1661 14653 1695
rect 14570 1647 14653 1661
rect 14502 1646 14653 1647
rect 14427 1627 14653 1646
rect 14427 1612 14604 1627
rect 14427 1611 14536 1612
rect 14427 1577 14468 1611
rect 14502 1578 14536 1611
rect 14570 1593 14604 1612
rect 14638 1593 14653 1627
rect 14570 1578 14653 1593
rect 14502 1577 14653 1578
rect 14427 1559 14653 1577
rect 14427 1552 14604 1559
rect 482 1551 682 1552
rect 482 1517 497 1551
rect 531 1541 682 1551
rect 531 1517 565 1541
rect 482 1507 565 1517
rect 599 1507 633 1541
rect 667 1507 682 1541
rect 482 1483 682 1507
rect 482 1449 497 1483
rect 531 1472 682 1483
rect 531 1449 565 1472
rect 482 1438 565 1449
rect 599 1438 633 1472
rect 667 1438 682 1472
rect 482 1415 682 1438
rect 482 1381 497 1415
rect 531 1403 682 1415
rect 531 1381 565 1403
rect 482 1369 565 1381
rect 599 1369 633 1403
rect 667 1369 682 1403
rect 14453 1543 14604 1552
rect 14453 1542 14536 1543
rect 14453 1508 14468 1542
rect 14502 1509 14536 1542
rect 14570 1525 14604 1543
rect 14638 1525 14653 1559
rect 14570 1509 14653 1525
rect 14502 1508 14653 1509
rect 14453 1491 14653 1508
rect 14453 1474 14604 1491
rect 14453 1473 14536 1474
rect 14453 1439 14468 1473
rect 14502 1440 14536 1473
rect 14570 1457 14604 1474
rect 14638 1457 14653 1491
rect 14570 1440 14653 1457
rect 14502 1439 14653 1440
rect 14453 1423 14653 1439
rect 14453 1405 14604 1423
rect 14453 1404 14536 1405
rect 482 1347 682 1369
rect 482 1313 497 1347
rect 531 1334 682 1347
rect 531 1313 565 1334
rect 482 1300 565 1313
rect 599 1300 633 1334
rect 667 1300 682 1334
rect 482 1279 682 1300
rect 482 1245 497 1279
rect 531 1265 682 1279
rect 531 1245 565 1265
rect 482 1231 565 1245
rect 599 1231 633 1265
rect 667 1231 682 1265
rect 482 1211 682 1231
rect 482 1177 497 1211
rect 531 1196 682 1211
rect 531 1177 565 1196
rect 482 1162 565 1177
rect 599 1162 633 1196
rect 667 1162 682 1196
rect 482 1143 682 1162
rect 482 1109 497 1143
rect 531 1127 682 1143
rect 531 1109 565 1127
rect 482 1093 565 1109
rect 599 1093 633 1127
rect 667 1093 682 1127
rect 482 1075 682 1093
rect 482 1041 497 1075
rect 531 1058 682 1075
rect 531 1041 565 1058
rect 482 1024 565 1041
rect 599 1024 633 1058
rect 667 1024 682 1058
rect 482 1007 682 1024
rect 482 973 497 1007
rect 531 989 682 1007
rect 531 973 565 989
rect 482 955 565 973
rect 599 955 633 989
rect 667 955 682 989
rect 482 939 682 955
rect 482 769 497 939
rect 531 920 682 939
rect 667 867 682 920
rect 14453 1370 14468 1404
rect 14502 1371 14536 1404
rect 14570 1389 14604 1405
rect 14638 1389 14653 1423
rect 14570 1371 14653 1389
rect 14502 1370 14653 1371
rect 14453 1355 14653 1370
rect 14453 1336 14604 1355
rect 14453 1335 14536 1336
rect 14453 1301 14468 1335
rect 14502 1302 14536 1335
rect 14570 1321 14604 1336
rect 14638 1321 14653 1355
rect 14570 1302 14653 1321
rect 14502 1301 14653 1302
rect 14453 1287 14653 1301
rect 14453 1267 14604 1287
rect 14453 1266 14536 1267
rect 14453 1232 14468 1266
rect 14502 1233 14536 1266
rect 14570 1253 14604 1267
rect 14638 1253 14653 1287
rect 14570 1233 14653 1253
rect 14502 1232 14653 1233
rect 14453 1218 14653 1232
rect 14453 1198 14604 1218
rect 14453 1197 14536 1198
rect 14453 1163 14468 1197
rect 14502 1164 14536 1197
rect 14570 1184 14604 1198
rect 14638 1184 14653 1218
rect 14570 1164 14653 1184
rect 14502 1163 14653 1164
rect 14453 1149 14653 1163
rect 14453 1129 14604 1149
rect 14453 1128 14536 1129
rect 14453 1094 14468 1128
rect 14502 1095 14536 1128
rect 14570 1115 14604 1129
rect 14638 1115 14653 1149
rect 14570 1095 14653 1115
rect 14502 1094 14653 1095
rect 14453 1080 14653 1094
rect 14453 1060 14604 1080
rect 14453 1059 14536 1060
rect 14453 1025 14468 1059
rect 14502 1026 14536 1059
rect 14570 1046 14604 1060
rect 14638 1046 14653 1080
rect 14570 1026 14653 1046
rect 14502 1025 14653 1026
rect 14453 1011 14653 1025
rect 14453 991 14604 1011
rect 14453 990 14536 991
rect 14453 956 14468 990
rect 14502 957 14536 990
rect 14570 977 14604 991
rect 14638 977 14653 1011
rect 14570 957 14653 977
rect 14502 956 14653 957
rect 14453 942 14653 956
rect 14453 922 14604 942
rect 14453 921 14536 922
rect 14453 887 14468 921
rect 14502 888 14536 921
rect 14570 908 14604 922
rect 14638 908 14653 942
rect 14570 888 14653 908
rect 14502 887 14653 888
rect 14453 873 14653 887
rect 14453 867 14604 873
rect 667 853 14604 867
rect 667 852 14536 853
rect 667 818 702 852
rect 736 818 771 852
rect 805 818 840 852
rect 874 818 909 852
rect 943 818 978 852
rect 1012 818 1047 852
rect 1081 818 1116 852
rect 1150 818 1185 852
rect 1219 818 1254 852
rect 1288 818 1323 852
rect 1357 818 1392 852
rect 1426 818 1461 852
rect 1495 818 1530 852
rect 1564 818 1599 852
rect 1633 818 1668 852
rect 1702 818 1737 852
rect 1771 818 1806 852
rect 1840 818 1875 852
rect 1909 818 1944 852
rect 1978 818 2013 852
rect 2047 818 2082 852
rect 2116 818 2151 852
rect 2185 818 2220 852
rect 2254 818 2289 852
rect 2323 818 2358 852
rect 2392 818 2427 852
rect 2461 818 2496 852
rect 2530 818 2565 852
rect 2599 818 2634 852
rect 2668 818 2703 852
rect 2737 818 2772 852
rect 599 784 2772 818
rect 14502 819 14536 852
rect 14570 839 14604 853
rect 14638 839 14653 873
rect 14570 819 14653 839
rect 14502 804 14653 819
rect 14502 784 14604 804
rect 482 750 565 769
rect 599 750 634 784
rect 668 750 703 784
rect 737 750 772 784
rect 806 750 841 784
rect 875 750 910 784
rect 944 750 979 784
rect 1013 750 1048 784
rect 1082 750 1117 784
rect 1151 750 1186 784
rect 1220 750 1255 784
rect 1289 750 1324 784
rect 1358 750 1393 784
rect 1427 750 1462 784
rect 1496 750 1531 784
rect 1565 750 1600 784
rect 1634 750 1669 784
rect 1703 750 1738 784
rect 1772 750 1807 784
rect 1841 750 1876 784
rect 1910 750 1945 784
rect 1979 750 2014 784
rect 2048 750 2083 784
rect 2117 750 2152 784
rect 2186 750 2221 784
rect 2255 750 2290 784
rect 2324 750 2359 784
rect 2393 750 2428 784
rect 2462 750 2497 784
rect 2531 750 2566 784
rect 2600 750 2635 784
rect 2669 750 2704 784
rect 2738 750 2772 784
rect 14570 770 14604 784
rect 14638 770 14653 804
rect 14570 750 14653 770
rect 482 716 4725 750
rect 482 682 516 716
rect 550 682 585 716
rect 619 682 654 716
rect 688 682 723 716
rect 757 682 792 716
rect 826 682 861 716
rect 895 682 930 716
rect 964 682 999 716
rect 1033 682 1068 716
rect 1102 682 1137 716
rect 1171 682 1206 716
rect 1240 682 1275 716
rect 1309 682 1344 716
rect 1378 682 1413 716
rect 1447 682 1482 716
rect 1516 682 1551 716
rect 1585 682 1620 716
rect 1654 682 1689 716
rect 1723 682 1758 716
rect 1792 682 1827 716
rect 1861 682 1896 716
rect 1930 682 1965 716
rect 1999 682 2034 716
rect 2068 682 2103 716
rect 2137 682 2172 716
rect 2206 682 2241 716
rect 2275 682 2310 716
rect 2344 682 2379 716
rect 2413 682 2448 716
rect 2482 682 2517 716
rect 2551 682 2586 716
rect 2620 682 2655 716
rect 2689 682 2724 716
rect 2758 682 2793 716
rect 2827 682 2862 716
rect 2896 682 2931 716
rect 2965 682 3000 716
rect 3034 682 3069 716
rect 3103 682 3138 716
rect 3172 682 3207 716
rect 3241 682 3276 716
rect 3310 682 3345 716
rect 3379 682 3414 716
rect 3448 682 3483 716
rect 3517 682 3552 716
rect 3586 682 3621 716
rect 3655 682 3690 716
rect 3724 682 3759 716
rect 3793 682 3828 716
rect 3862 682 3897 716
rect 3931 682 3966 716
rect 4000 682 4035 716
rect 4069 682 4104 716
rect 4138 682 4173 716
rect 4207 682 4242 716
rect 4276 682 4311 716
rect 4345 682 4380 716
rect 4414 682 4449 716
rect 4483 682 4518 716
rect 4552 682 4587 716
rect 4621 682 4656 716
rect 4690 682 4725 716
rect 14551 735 14653 750
rect 14551 701 14604 735
rect 14638 701 14653 735
rect 14551 682 14653 701
rect 482 667 14653 682
<< mvpsubdiffcont >>
rect 51 5015 85 5049
rect 142 5034 176 5068
rect 214 5034 248 5068
rect 286 5034 320 5068
rect 358 5034 392 5068
rect 430 5034 464 5068
rect 502 5034 536 5068
rect 574 5034 608 5068
rect 646 5034 680 5068
rect 718 5034 752 5068
rect 790 5034 824 5068
rect 862 5034 896 5068
rect 934 5034 968 5068
rect 1006 5034 1040 5068
rect 1078 5034 1112 5068
rect 1150 5034 1184 5068
rect 1222 5034 1256 5068
rect 1294 5034 1328 5068
rect 1366 5034 1400 5068
rect 1438 5034 1472 5068
rect 1510 5034 1544 5068
rect 1582 5034 1616 5068
rect 1654 5034 1688 5068
rect 1726 5034 1760 5068
rect 1798 5034 1832 5068
rect 1870 5034 1904 5068
rect 1942 5034 1976 5068
rect 2014 5034 2048 5068
rect 2086 5034 2120 5068
rect 2158 5034 2192 5068
rect 2230 5034 2264 5068
rect 2302 5034 2336 5068
rect 2374 5034 2408 5068
rect 2446 5034 2480 5068
rect 2518 5034 2552 5068
rect 2590 5034 2624 5068
rect 2662 5034 2696 5068
rect 2734 5034 2768 5068
rect 2806 5034 2840 5068
rect 2878 5034 2912 5068
rect 2950 5034 2984 5068
rect 3022 5034 3056 5068
rect 3094 5034 3128 5068
rect 3166 5034 3200 5068
rect 3238 5034 3272 5068
rect 3310 5034 3344 5068
rect 3382 5034 3416 5068
rect 3454 5034 3488 5068
rect 3526 5034 3560 5068
rect 3598 5034 3632 5068
rect 3670 5034 3704 5068
rect 3742 5034 3776 5068
rect 3814 5034 3848 5068
rect 3886 5034 3920 5068
rect 3958 5034 3992 5068
rect 4030 5034 4064 5068
rect 4102 5034 4136 5068
rect 4174 5034 4208 5068
rect 4246 5034 4280 5068
rect 4318 5034 4352 5068
rect 4390 5034 4424 5068
rect 4462 5034 4496 5068
rect 4534 5034 4568 5068
rect 4606 5034 4640 5068
rect 4678 5034 4712 5068
rect 4750 5034 4784 5068
rect 4822 5034 4856 5068
rect 4894 5034 4928 5068
rect 4966 5034 5000 5068
rect 5038 5034 5072 5068
rect 5110 5034 5144 5068
rect 5182 5034 5216 5068
rect 5254 5034 5288 5068
rect 5326 5034 5360 5068
rect 5398 5034 5432 5068
rect 5470 5034 5504 5068
rect 5542 5034 5576 5068
rect 5614 5034 5648 5068
rect 5686 5034 5720 5068
rect 5758 5034 5792 5068
rect 5830 5034 5864 5068
rect 5902 5034 5936 5068
rect 5974 5034 6008 5068
rect 6046 5034 6080 5068
rect 6118 5034 6152 5068
rect 6190 5034 6224 5068
rect 6262 5034 6296 5068
rect 6334 5034 6368 5068
rect 6406 5034 6440 5068
rect 6478 5034 6512 5068
rect 6550 5034 6584 5068
rect 6622 5034 6656 5068
rect 6694 5034 6728 5068
rect 6766 5034 6800 5068
rect 6838 5034 6872 5068
rect 6910 5034 6944 5068
rect 6982 5034 7016 5068
rect 7054 5034 7088 5068
rect 7126 5034 7160 5068
rect 7198 5034 7232 5068
rect 7270 5034 7304 5068
rect 7342 5034 7376 5068
rect 7414 5034 7448 5068
rect 7486 5034 7520 5068
rect 7558 5034 7592 5068
rect 7630 5034 7664 5068
rect 7702 5034 7736 5068
rect 7774 5034 7808 5068
rect 7846 5034 7880 5068
rect 7918 5034 7952 5068
rect 7990 5034 8024 5068
rect 8062 5034 8096 5068
rect 8134 5034 8168 5068
rect 8206 5034 8240 5068
rect 8278 5034 8312 5068
rect 8350 5034 8384 5068
rect 8422 5034 8456 5068
rect 8494 5034 8528 5068
rect 8566 5034 8600 5068
rect 8638 5034 8672 5068
rect 8710 5034 8744 5068
rect 8782 5034 8816 5068
rect 8854 5034 8888 5068
rect 8926 5034 8960 5068
rect 8998 5034 9032 5068
rect 9070 5034 9104 5068
rect 9142 5034 9176 5068
rect 9214 5034 9248 5068
rect 9286 5034 9320 5068
rect 9358 5034 9392 5068
rect 9430 5034 9464 5068
rect 9502 5034 9536 5068
rect 9574 5034 9608 5068
rect 9646 5034 9680 5068
rect 9718 5034 9752 5068
rect 9790 5034 9824 5068
rect 9862 5034 9896 5068
rect 9934 5034 9968 5068
rect 10006 5034 10040 5068
rect 10078 5034 10112 5068
rect 10151 5034 10185 5068
rect 10224 5034 10258 5068
rect 10297 5034 10331 5068
rect 10370 5034 10404 5068
rect 10443 5034 10477 5068
rect 10516 5034 10550 5068
rect 10589 5034 10623 5068
rect 10662 5034 10696 5068
rect 10735 5034 10769 5068
rect 10808 5034 10842 5068
rect 10881 5034 10915 5068
rect 10954 5034 10988 5068
rect 11027 5034 11061 5068
rect 11100 5034 11134 5068
rect 11173 5034 11207 5068
rect 11246 5034 11280 5068
rect 11319 5034 11353 5068
rect 11392 5034 11426 5068
rect 11465 5034 11499 5068
rect 11538 5034 11572 5068
rect 11611 5034 11645 5068
rect 11684 5034 11718 5068
rect 11757 5034 11791 5068
rect 11830 5034 11864 5068
rect 11903 5034 11937 5068
rect 11976 5034 12010 5068
rect 12049 5034 12083 5068
rect 12122 5034 12156 5068
rect 12195 5034 12229 5068
rect 12268 5034 12302 5068
rect 12341 5034 12375 5068
rect 12414 5034 12448 5068
rect 12487 5034 12521 5068
rect 12560 5034 12594 5068
rect 12633 5034 12667 5068
rect 12706 5034 12740 5068
rect 12779 5034 12813 5068
rect 12852 5034 12886 5068
rect 12925 5034 12959 5068
rect 12998 5034 13032 5068
rect 13071 5034 13105 5068
rect 13144 5034 13178 5068
rect 13217 5034 13251 5068
rect 13290 5034 13324 5068
rect 13363 5034 13397 5068
rect 13436 5034 13470 5068
rect 13509 5034 13543 5068
rect 13582 5034 13616 5068
rect 13655 5034 13689 5068
rect 13728 5034 13762 5068
rect 13801 5034 13835 5068
rect 13874 5034 13908 5068
rect 13947 5034 13981 5068
rect 14020 5034 14054 5068
rect 14093 5034 14127 5068
rect 14166 5034 14200 5068
rect 14239 5034 14273 5068
rect 14312 5034 14346 5068
rect 14385 5034 14419 5068
rect 14458 5034 14492 5068
rect 14531 5034 14565 5068
rect 14604 5034 14638 5068
rect 14677 5034 14711 5068
rect 14750 5034 14784 5068
rect 14823 5034 14857 5068
rect 51 4942 85 4976
rect 119 4966 153 5000
rect 191 4966 225 5000
rect 263 4966 297 5000
rect 335 4966 369 5000
rect 407 4966 441 5000
rect 479 4966 513 5000
rect 551 4966 585 5000
rect 623 4966 657 5000
rect 695 4966 729 5000
rect 767 4966 801 5000
rect 839 4966 873 5000
rect 911 4966 945 5000
rect 983 4966 1017 5000
rect 1055 4966 1089 5000
rect 1127 4966 1161 5000
rect 1199 4966 1233 5000
rect 1271 4966 1305 5000
rect 1343 4966 1377 5000
rect 1415 4966 1449 5000
rect 1487 4966 1521 5000
rect 1559 4966 1593 5000
rect 1631 4966 1665 5000
rect 1703 4966 1737 5000
rect 1775 4966 1809 5000
rect 1847 4966 1881 5000
rect 1919 4966 1953 5000
rect 1991 4966 2025 5000
rect 2063 4966 2097 5000
rect 2135 4966 2169 5000
rect 2207 4966 2241 5000
rect 2279 4966 2313 5000
rect 2351 4966 2385 5000
rect 2423 4966 2457 5000
rect 2495 4966 2529 5000
rect 2567 4966 2601 5000
rect 2639 4966 2673 5000
rect 2711 4966 2745 5000
rect 2783 4966 2817 5000
rect 2855 4966 2889 5000
rect 2927 4966 2961 5000
rect 2999 4966 3033 5000
rect 3071 4966 3105 5000
rect 3143 4966 3177 5000
rect 3215 4966 3249 5000
rect 3287 4966 3321 5000
rect 3359 4966 3393 5000
rect 3431 4966 3465 5000
rect 3503 4966 3537 5000
rect 3575 4966 3609 5000
rect 3647 4966 3681 5000
rect 3719 4966 3753 5000
rect 3791 4966 3825 5000
rect 3863 4966 3897 5000
rect 3935 4966 3969 5000
rect 4007 4966 4041 5000
rect 4079 4966 4113 5000
rect 4151 4966 4185 5000
rect 4223 4966 4257 5000
rect 4295 4966 4329 5000
rect 4367 4966 4401 5000
rect 4439 4966 4473 5000
rect 4511 4966 4545 5000
rect 4583 4966 4617 5000
rect 4655 4966 4689 5000
rect 4727 4966 4761 5000
rect 4799 4966 4833 5000
rect 4871 4966 4905 5000
rect 4943 4966 4977 5000
rect 5015 4966 5049 5000
rect 5087 4966 5121 5000
rect 5159 4966 5193 5000
rect 5231 4966 5265 5000
rect 5303 4966 5337 5000
rect 5375 4966 5409 5000
rect 5447 4966 5481 5000
rect 5519 4966 5553 5000
rect 5591 4966 5625 5000
rect 5663 4966 5697 5000
rect 5735 4966 5769 5000
rect 5807 4966 5841 5000
rect 5879 4966 5913 5000
rect 5951 4966 5985 5000
rect 6023 4966 6057 5000
rect 6095 4966 6129 5000
rect 6167 4966 6201 5000
rect 6239 4966 6273 5000
rect 6311 4966 6345 5000
rect 6383 4966 6417 5000
rect 6455 4966 6489 5000
rect 6527 4966 6561 5000
rect 6599 4966 6633 5000
rect 6671 4966 6705 5000
rect 6743 4966 6777 5000
rect 6815 4966 6849 5000
rect 6887 4966 6921 5000
rect 6959 4966 6993 5000
rect 7031 4966 7065 5000
rect 7103 4966 7137 5000
rect 7175 4966 7209 5000
rect 7247 4966 7281 5000
rect 7319 4966 7353 5000
rect 7391 4966 7425 5000
rect 7463 4966 7497 5000
rect 7535 4966 7569 5000
rect 7607 4966 7641 5000
rect 7679 4966 7713 5000
rect 7751 4966 7785 5000
rect 7823 4966 7857 5000
rect 7895 4966 7929 5000
rect 7967 4966 8001 5000
rect 8039 4966 8073 5000
rect 8111 4966 8145 5000
rect 8183 4966 8217 5000
rect 8255 4966 8289 5000
rect 8327 4966 8361 5000
rect 8399 4966 8433 5000
rect 8471 4966 8505 5000
rect 8543 4966 8577 5000
rect 8615 4966 8649 5000
rect 8687 4966 8721 5000
rect 8759 4966 8793 5000
rect 8831 4966 8865 5000
rect 8903 4966 8937 5000
rect 8975 4966 9009 5000
rect 9047 4966 9081 5000
rect 9119 4966 9153 5000
rect 9191 4966 9225 5000
rect 9263 4966 9297 5000
rect 9335 4966 9369 5000
rect 9407 4966 9441 5000
rect 9479 4966 9513 5000
rect 9551 4966 9585 5000
rect 9623 4966 9657 5000
rect 9695 4966 9729 5000
rect 9767 4966 9801 5000
rect 9839 4966 9873 5000
rect 9911 4966 9945 5000
rect 9983 4966 10017 5000
rect 10055 4966 10089 5000
rect 10127 4966 10161 5000
rect 10199 4966 10233 5000
rect 10271 4966 10305 5000
rect 10343 4966 10377 5000
rect 10415 4966 10449 5000
rect 10487 4966 10521 5000
rect 10559 4966 10593 5000
rect 10631 4966 10665 5000
rect 10703 4966 10737 5000
rect 10775 4966 10809 5000
rect 10847 4966 10881 5000
rect 10919 4966 10953 5000
rect 10991 4966 11025 5000
rect 11063 4966 11097 5000
rect 11135 4966 11169 5000
rect 11207 4966 11241 5000
rect 11279 4966 11313 5000
rect 11351 4966 11385 5000
rect 11423 4966 11457 5000
rect 11495 4966 11529 5000
rect 11567 4966 11601 5000
rect 11639 4966 11673 5000
rect 11711 4966 11745 5000
rect 11783 4966 11817 5000
rect 11855 4966 11889 5000
rect 11927 4966 11961 5000
rect 11999 4966 12033 5000
rect 12071 4966 12105 5000
rect 12143 4966 12177 5000
rect 12215 4966 12249 5000
rect 12287 4966 12321 5000
rect 12359 4966 12393 5000
rect 12431 4966 12465 5000
rect 12503 4966 12537 5000
rect 12575 4966 12609 5000
rect 12647 4966 12681 5000
rect 12719 4966 12753 5000
rect 12791 4966 12825 5000
rect 12863 4966 12897 5000
rect 12935 4966 12969 5000
rect 13007 4966 13041 5000
rect 13079 4966 13113 5000
rect 13151 4966 13185 5000
rect 13223 4966 13257 5000
rect 13295 4966 13329 5000
rect 13367 4966 13401 5000
rect 13439 4966 13473 5000
rect 13511 4966 13545 5000
rect 13583 4966 13617 5000
rect 13655 4966 13689 5000
rect 13728 4966 13762 5000
rect 13801 4966 13835 5000
rect 13874 4966 13908 5000
rect 13947 4966 13981 5000
rect 14020 4966 14054 5000
rect 14093 4966 14127 5000
rect 14166 4966 14200 5000
rect 14239 4966 14273 5000
rect 14312 4966 14346 5000
rect 14385 4966 14419 5000
rect 14458 4966 14492 5000
rect 14531 4966 14565 5000
rect 14604 4966 14638 5000
rect 14677 4966 14711 5000
rect 14750 4966 14784 5000
rect 14823 4966 14857 5000
rect 14915 4983 14949 5017
rect 14983 4983 15017 5017
rect 15051 4983 15085 5017
rect 51 4869 85 4903
rect 119 4892 153 4926
rect 187 4898 221 4932
rect 259 4898 293 4932
rect 331 4898 365 4932
rect 403 4898 437 4932
rect 475 4898 509 4932
rect 547 4898 581 4932
rect 619 4898 653 4932
rect 691 4898 725 4932
rect 763 4898 797 4932
rect 835 4898 869 4932
rect 907 4898 941 4932
rect 979 4898 1013 4932
rect 1051 4898 1085 4932
rect 1123 4898 1157 4932
rect 1195 4898 1229 4932
rect 1267 4898 1301 4932
rect 1339 4898 1373 4932
rect 1411 4898 1445 4932
rect 1483 4898 1517 4932
rect 1555 4898 1589 4932
rect 1627 4898 1661 4932
rect 1699 4898 1733 4932
rect 1771 4898 1805 4932
rect 1843 4898 1877 4932
rect 1915 4898 1949 4932
rect 1987 4898 2021 4932
rect 2059 4898 2093 4932
rect 2131 4898 2165 4932
rect 2203 4898 2237 4932
rect 2275 4898 2309 4932
rect 2347 4898 2381 4932
rect 2419 4898 2453 4932
rect 2491 4898 2525 4932
rect 2563 4898 2597 4932
rect 2635 4898 2669 4932
rect 2707 4898 2741 4932
rect 2779 4898 2813 4932
rect 2851 4898 2885 4932
rect 2923 4898 2957 4932
rect 2995 4898 3029 4932
rect 3067 4898 3101 4932
rect 3139 4898 3173 4932
rect 3211 4898 3245 4932
rect 3283 4898 3317 4932
rect 3355 4898 3389 4932
rect 3427 4898 3461 4932
rect 3499 4898 3533 4932
rect 3571 4898 3605 4932
rect 3643 4898 3677 4932
rect 3715 4898 3749 4932
rect 3787 4898 3821 4932
rect 3859 4898 3893 4932
rect 3931 4898 3965 4932
rect 4003 4898 4037 4932
rect 4075 4898 4109 4932
rect 4147 4898 4181 4932
rect 4219 4898 4253 4932
rect 4291 4898 4325 4932
rect 4363 4898 4397 4932
rect 4435 4898 4469 4932
rect 4507 4898 4541 4932
rect 4579 4898 4613 4932
rect 4651 4898 4685 4932
rect 4723 4898 4757 4932
rect 4795 4898 4829 4932
rect 4867 4898 4901 4932
rect 4939 4898 4973 4932
rect 5011 4898 5045 4932
rect 5083 4898 5117 4932
rect 5155 4898 5189 4932
rect 5227 4898 5261 4932
rect 5299 4898 5333 4932
rect 5371 4898 5405 4932
rect 5443 4898 5477 4932
rect 5515 4898 5549 4932
rect 5587 4898 5621 4932
rect 5659 4898 5693 4932
rect 5731 4898 5765 4932
rect 5803 4898 5837 4932
rect 5875 4898 5909 4932
rect 5947 4898 5981 4932
rect 6019 4898 6053 4932
rect 6091 4898 6125 4932
rect 6163 4898 6197 4932
rect 6235 4898 6269 4932
rect 6307 4898 6341 4932
rect 6379 4898 6413 4932
rect 6451 4898 6485 4932
rect 6523 4898 6557 4932
rect 6595 4898 6629 4932
rect 6667 4898 6701 4932
rect 6739 4898 6773 4932
rect 6811 4898 6845 4932
rect 6883 4898 6917 4932
rect 6955 4898 6989 4932
rect 7027 4898 7061 4932
rect 7099 4898 7133 4932
rect 7171 4898 7205 4932
rect 7243 4898 7277 4932
rect 7315 4898 7349 4932
rect 7387 4898 7421 4932
rect 7459 4898 7493 4932
rect 7531 4898 7565 4932
rect 7603 4898 7637 4932
rect 7675 4898 7709 4932
rect 7747 4898 7781 4932
rect 7819 4898 7853 4932
rect 7891 4898 7925 4932
rect 7963 4898 7997 4932
rect 8035 4898 8069 4932
rect 8107 4898 8141 4932
rect 8179 4898 8213 4932
rect 8251 4898 8285 4932
rect 8323 4898 8357 4932
rect 8395 4898 8429 4932
rect 8467 4898 8501 4932
rect 8539 4898 8573 4932
rect 8611 4898 8645 4932
rect 8683 4898 8717 4932
rect 8755 4898 8789 4932
rect 8827 4898 8861 4932
rect 8899 4898 8933 4932
rect 8971 4898 9005 4932
rect 9043 4898 9077 4932
rect 9115 4898 9149 4932
rect 9187 4898 9221 4932
rect 9259 4898 9293 4932
rect 9331 4898 9365 4932
rect 9403 4898 9437 4932
rect 9475 4898 9509 4932
rect 9547 4898 9581 4932
rect 9619 4898 9653 4932
rect 9691 4898 9725 4932
rect 9763 4898 9797 4932
rect 9835 4898 9869 4932
rect 9907 4898 9941 4932
rect 9979 4898 10013 4932
rect 10051 4898 10085 4932
rect 10123 4898 10157 4932
rect 10195 4898 10229 4932
rect 10267 4898 10301 4932
rect 10339 4898 10373 4932
rect 10411 4898 10445 4932
rect 10483 4898 10517 4932
rect 10555 4898 10589 4932
rect 10627 4898 10661 4932
rect 10699 4898 10733 4932
rect 10771 4898 10805 4932
rect 10843 4898 10877 4932
rect 10915 4898 10949 4932
rect 10987 4898 11021 4932
rect 11059 4898 11093 4932
rect 11131 4898 11165 4932
rect 11203 4898 11237 4932
rect 11275 4898 11309 4932
rect 11347 4898 11381 4932
rect 11419 4898 11453 4932
rect 11491 4898 11525 4932
rect 11563 4898 11597 4932
rect 11635 4898 11669 4932
rect 11707 4898 11741 4932
rect 11779 4898 11813 4932
rect 11851 4898 11885 4932
rect 11923 4898 11957 4932
rect 11995 4898 12029 4932
rect 12067 4898 12101 4932
rect 12139 4898 12173 4932
rect 12211 4898 12245 4932
rect 12283 4898 12317 4932
rect 12355 4898 12389 4932
rect 12427 4898 12461 4932
rect 12499 4898 12533 4932
rect 12571 4898 12605 4932
rect 12643 4898 12677 4932
rect 12715 4898 12749 4932
rect 12787 4898 12821 4932
rect 12859 4898 12893 4932
rect 12931 4898 12965 4932
rect 13003 4898 13037 4932
rect 13075 4898 13109 4932
rect 13147 4898 13181 4932
rect 13219 4898 13253 4932
rect 13291 4898 13325 4932
rect 13363 4898 13397 4932
rect 13436 4898 13470 4932
rect 13509 4898 13543 4932
rect 13582 4898 13616 4932
rect 13655 4898 13689 4932
rect 13728 4898 13762 4932
rect 13801 4898 13835 4932
rect 13874 4898 13908 4932
rect 13947 4898 13981 4932
rect 14020 4898 14054 4932
rect 14093 4898 14127 4932
rect 14166 4898 14200 4932
rect 14239 4898 14273 4932
rect 14312 4898 14346 4932
rect 14385 4898 14419 4932
rect 14458 4898 14492 4932
rect 14531 4898 14565 4932
rect 14604 4898 14638 4932
rect 14677 4898 14711 4932
rect 14750 4898 14784 4932
rect 14823 4898 14857 4932
rect 14915 4911 14949 4945
rect 14983 4911 15017 4945
rect 15051 4911 15085 4945
rect 51 4796 85 4830
rect 119 4818 153 4852
rect 187 4823 221 4857
rect 262 4825 296 4859
rect 51 4723 85 4757
rect 119 4744 153 4778
rect 187 4748 221 4782
rect 262 4757 296 4791
rect 51 4650 85 4684
rect 119 4670 153 4704
rect 187 4673 221 4707
rect 262 4689 296 4723
rect 51 4577 85 4611
rect 119 4596 153 4630
rect 187 4598 221 4632
rect 262 4621 296 4655
rect 14840 4825 14874 4859
rect 14915 4839 14949 4873
rect 14983 4839 15017 4873
rect 15051 4839 15085 4873
rect 14840 4757 14874 4791
rect 14915 4767 14949 4801
rect 14983 4767 15017 4801
rect 15051 4767 15085 4801
rect 14840 4689 14874 4723
rect 14915 4695 14949 4729
rect 14983 4695 15017 4729
rect 15051 4695 15085 4729
rect 51 4504 85 4538
rect 119 4522 153 4556
rect 187 4523 221 4557
rect 262 4553 296 4587
rect 262 4485 296 4519
rect 51 4431 85 4465
rect 119 4448 153 4482
rect 187 4449 221 4483
rect 262 4417 296 4451
rect 51 4359 85 4393
rect 119 4374 153 4408
rect 187 4375 221 4409
rect 262 4349 296 4383
rect 51 4287 85 4321
rect 119 4300 153 4334
rect 187 4301 221 4335
rect 262 4281 296 4315
rect 51 4215 85 4249
rect 119 4226 153 4260
rect 187 4227 221 4261
rect 262 4213 296 4247
rect 51 4143 85 4177
rect 119 4152 153 4186
rect 187 4153 221 4187
rect 262 4145 296 4179
rect 51 4071 85 4105
rect 119 4078 153 4112
rect 187 4079 221 4113
rect 262 4077 296 4111
rect 51 3999 85 4033
rect 119 4004 153 4038
rect 187 4005 221 4039
rect 262 4009 296 4043
rect 51 3927 85 3961
rect 119 3930 153 3964
rect 187 3931 221 3965
rect 262 3941 296 3975
rect 51 3855 85 3889
rect 119 3856 153 3890
rect 187 3857 221 3891
rect 262 3873 296 3907
rect 51 3783 85 3817
rect 119 3783 153 3817
rect 187 3783 221 3817
rect 262 3805 296 3839
rect 262 3737 296 3771
rect 51 3673 85 3707
rect 119 3673 153 3707
rect 187 3673 221 3707
rect 262 3669 296 3703
rect 51 3600 85 3634
rect 119 3600 153 3634
rect 187 3600 221 3634
rect 262 3601 296 3635
rect 51 3528 85 3562
rect 119 3528 153 3562
rect 187 3528 221 3562
rect 262 3533 296 3567
rect 51 3456 85 3490
rect 119 3456 153 3490
rect 187 3456 221 3490
rect 262 3465 296 3499
rect 51 3384 85 3418
rect 119 3384 153 3418
rect 187 3384 221 3418
rect 262 3397 296 3431
rect 51 3312 85 3346
rect 119 3312 153 3346
rect 187 3312 221 3346
rect 262 3329 296 3363
rect 51 3240 85 3274
rect 119 3240 153 3274
rect 187 3240 221 3274
rect 262 3261 296 3295
rect 51 3168 85 3202
rect 119 3168 153 3202
rect 187 3168 221 3202
rect 262 3193 296 3227
rect 51 3096 85 3130
rect 119 3096 153 3130
rect 187 3096 221 3130
rect 262 3125 296 3159
rect 51 3024 85 3058
rect 119 3024 153 3058
rect 187 3024 221 3058
rect 262 3057 296 3091
rect 262 2989 296 3023
rect 51 2952 85 2986
rect 119 2952 153 2986
rect 187 2952 221 2986
rect 262 2921 296 2955
rect 51 2880 85 2914
rect 119 2880 153 2914
rect 187 2880 221 2914
rect 262 2853 296 2887
rect 51 2808 85 2842
rect 119 2808 153 2842
rect 187 2808 221 2842
rect 262 2785 296 2819
rect 51 2736 85 2770
rect 119 2736 153 2770
rect 187 2736 221 2770
rect 262 2717 296 2751
rect 51 2664 85 2698
rect 119 2664 153 2698
rect 187 2664 221 2698
rect 262 2649 296 2683
rect 51 2592 85 2626
rect 119 2592 153 2626
rect 187 2592 221 2626
rect 262 2581 296 2615
rect 51 2520 85 2554
rect 119 2520 153 2554
rect 187 2520 221 2554
rect 262 2513 296 2547
rect 51 2448 85 2482
rect 119 2448 153 2482
rect 187 2448 221 2482
rect 262 2445 296 2479
rect 51 2376 85 2410
rect 119 2376 153 2410
rect 187 2376 221 2410
rect 262 2377 296 2411
rect 51 2304 85 2338
rect 119 2304 153 2338
rect 187 2304 221 2338
rect 262 2309 296 2343
rect 51 2232 85 2266
rect 119 2232 153 2266
rect 187 2232 221 2266
rect 262 2241 296 2275
rect 51 2160 85 2194
rect 119 2160 153 2194
rect 187 2160 221 2194
rect 262 2173 296 2207
rect 51 2088 85 2122
rect 119 2088 153 2122
rect 187 2088 221 2122
rect 262 2105 296 2139
rect 51 2016 85 2050
rect 119 2016 153 2050
rect 187 2016 221 2050
rect 262 2037 296 2071
rect 51 1944 85 1978
rect 119 1944 153 1978
rect 187 1944 221 1978
rect 262 1969 296 2003
rect 51 1872 85 1906
rect 119 1872 153 1906
rect 187 1872 221 1906
rect 262 1901 296 1935
rect 51 1800 85 1834
rect 119 1800 153 1834
rect 187 1800 221 1834
rect 262 1833 296 1867
rect 262 1765 296 1799
rect 51 1728 85 1762
rect 119 1728 153 1762
rect 187 1728 221 1762
rect 262 1697 296 1731
rect 51 1656 85 1690
rect 119 1656 153 1690
rect 187 1656 221 1690
rect 262 1629 296 1663
rect 51 1584 85 1618
rect 119 1584 153 1618
rect 187 1584 221 1618
rect 262 1561 296 1595
rect 51 1512 85 1546
rect 119 1512 153 1546
rect 187 1512 221 1546
rect 262 1493 296 1527
rect 51 1440 85 1474
rect 119 1440 153 1474
rect 187 1440 221 1474
rect 262 1425 296 1459
rect 51 1368 85 1402
rect 119 1368 153 1402
rect 187 1368 221 1402
rect 262 1357 296 1391
rect 51 1296 85 1330
rect 119 1296 153 1330
rect 187 1296 221 1330
rect 262 1289 296 1323
rect 51 1224 85 1258
rect 119 1224 153 1258
rect 187 1224 221 1258
rect 262 1221 296 1255
rect 51 1152 85 1186
rect 119 1152 153 1186
rect 187 1152 221 1186
rect 262 1153 296 1187
rect 51 1080 85 1114
rect 119 1080 153 1114
rect 187 1080 221 1114
rect 262 1085 296 1119
rect 51 1008 85 1042
rect 119 1008 153 1042
rect 187 1008 221 1042
rect 262 1017 296 1051
rect 51 936 85 970
rect 119 936 153 970
rect 187 936 221 970
rect 262 949 296 983
rect 51 864 85 898
rect 119 864 153 898
rect 187 864 221 898
rect 262 881 296 915
rect 51 792 85 826
rect 119 792 153 826
rect 187 792 221 826
rect 262 813 296 847
rect 51 720 85 754
rect 119 720 153 754
rect 187 720 221 754
rect 262 745 296 779
rect 51 648 85 682
rect 119 648 153 682
rect 187 648 221 682
rect 262 677 296 711
rect 14840 4621 14874 4655
rect 14915 4623 14949 4657
rect 14983 4623 15017 4657
rect 15051 4623 15085 4657
rect 14840 4553 14874 4587
rect 14915 4551 14949 4585
rect 14983 4551 15017 4585
rect 15051 4551 15085 4585
rect 14840 4485 14874 4519
rect 14915 4479 14949 4513
rect 14983 4479 15017 4513
rect 15051 4479 15085 4513
rect 14840 4417 14874 4451
rect 14915 4407 14949 4441
rect 14983 4407 15017 4441
rect 15051 4407 15085 4441
rect 14840 4349 14874 4383
rect 14915 4334 14949 4368
rect 14983 4335 15017 4369
rect 15051 4335 15085 4369
rect 14840 4281 14874 4315
rect 14915 4261 14949 4295
rect 14983 4263 15017 4297
rect 15051 4263 15085 4297
rect 14840 4213 14874 4247
rect 14915 4188 14949 4222
rect 14983 4191 15017 4225
rect 15051 4191 15085 4225
rect 14840 4145 14874 4179
rect 14915 4115 14949 4149
rect 14983 4119 15017 4153
rect 15051 4119 15085 4153
rect 14840 4077 14874 4111
rect 14840 4009 14874 4043
rect 14915 4042 14949 4076
rect 14983 4047 15017 4081
rect 15051 4047 15085 4081
rect 14840 3941 14874 3975
rect 14915 3969 14949 4003
rect 14983 3974 15017 4008
rect 15051 3975 15085 4009
rect 14840 3873 14874 3907
rect 14915 3896 14949 3930
rect 14983 3901 15017 3935
rect 15051 3903 15085 3937
rect 14840 3805 14874 3839
rect 14915 3823 14949 3857
rect 14983 3828 15017 3862
rect 15051 3831 15085 3865
rect 14840 3737 14874 3771
rect 14915 3750 14949 3784
rect 14983 3755 15017 3789
rect 15051 3759 15085 3793
rect 14840 3669 14874 3703
rect 14915 3677 14949 3711
rect 14983 3682 15017 3716
rect 15051 3687 15085 3721
rect 14840 3601 14874 3635
rect 14915 3604 14949 3638
rect 14983 3609 15017 3643
rect 15051 3615 15085 3649
rect 14840 3533 14874 3567
rect 14915 3531 14949 3565
rect 14983 3536 15017 3570
rect 15051 3543 15085 3577
rect 14840 3465 14874 3499
rect 14915 3458 14949 3492
rect 14983 3463 15017 3497
rect 15051 3471 15085 3505
rect 14840 3397 14874 3431
rect 14915 3385 14949 3419
rect 14983 3390 15017 3424
rect 15051 3399 15085 3433
rect 14840 3329 14874 3363
rect 14915 3312 14949 3346
rect 14983 3317 15017 3351
rect 15051 3327 15085 3361
rect 14840 3261 14874 3295
rect 14915 3239 14949 3273
rect 14983 3244 15017 3278
rect 15051 3255 15085 3289
rect 14840 3193 14874 3227
rect 14915 3166 14949 3200
rect 14983 3171 15017 3205
rect 15051 3183 15085 3217
rect 14840 3125 14874 3159
rect 14915 3093 14949 3127
rect 14983 3098 15017 3132
rect 15051 3111 15085 3145
rect 14840 3057 14874 3091
rect 14840 2989 14874 3023
rect 14915 3020 14949 3054
rect 14983 3025 15017 3059
rect 15051 3039 15085 3073
rect 14840 2921 14874 2955
rect 14915 2947 14949 2981
rect 14983 2952 15017 2986
rect 15051 2967 15085 3001
rect 14840 2853 14874 2887
rect 14915 2874 14949 2908
rect 14983 2879 15017 2913
rect 15051 2895 15085 2929
rect 14840 2785 14874 2819
rect 14915 2801 14949 2835
rect 14983 2806 15017 2840
rect 15051 2823 15085 2857
rect 14840 2717 14874 2751
rect 14915 2728 14949 2762
rect 14983 2733 15017 2767
rect 15051 2751 15085 2785
rect 14840 2649 14874 2683
rect 14915 2655 14949 2689
rect 14983 2660 15017 2694
rect 15051 2679 15085 2713
rect 14840 2581 14874 2615
rect 14915 2582 14949 2616
rect 14983 2587 15017 2621
rect 15051 2607 15085 2641
rect 14840 2513 14874 2547
rect 14915 2509 14949 2543
rect 14983 2514 15017 2548
rect 15051 2535 15085 2569
rect 14840 2445 14874 2479
rect 14915 2436 14949 2470
rect 14983 2441 15017 2475
rect 15051 2463 15085 2497
rect 14840 2377 14874 2411
rect 14915 2363 14949 2397
rect 14983 2368 15017 2402
rect 15051 2391 15085 2425
rect 14840 2309 14874 2343
rect 14915 2290 14949 2324
rect 14983 2295 15017 2329
rect 15051 2319 15085 2353
rect 14840 2241 14874 2275
rect 14915 2217 14949 2251
rect 14983 2222 15017 2256
rect 15051 2246 15085 2280
rect 14840 2173 14874 2207
rect 14915 2144 14949 2178
rect 14983 2149 15017 2183
rect 15051 2173 15085 2207
rect 14840 2105 14874 2139
rect 14915 2071 14949 2105
rect 14983 2076 15017 2110
rect 15051 2100 15085 2134
rect 14840 2037 14874 2071
rect 14840 1969 14874 2003
rect 14915 1998 14949 2032
rect 14983 2003 15017 2037
rect 15051 2027 15085 2061
rect 14840 1901 14874 1935
rect 14915 1925 14949 1959
rect 14983 1930 15017 1964
rect 15051 1954 15085 1988
rect 14840 1833 14874 1867
rect 14915 1852 14949 1886
rect 14983 1857 15017 1891
rect 15051 1881 15085 1915
rect 14840 1765 14874 1799
rect 14915 1779 14949 1813
rect 14983 1784 15017 1818
rect 15051 1808 15085 1842
rect 14840 1697 14874 1731
rect 14915 1706 14949 1740
rect 14983 1711 15017 1745
rect 15051 1735 15085 1769
rect 14840 1629 14874 1663
rect 14915 1633 14949 1667
rect 14983 1638 15017 1672
rect 15051 1662 15085 1696
rect 14840 1561 14874 1595
rect 14915 1560 14949 1594
rect 14983 1565 15017 1599
rect 15051 1589 15085 1623
rect 14840 1493 14874 1527
rect 14915 1487 14949 1521
rect 14983 1492 15017 1526
rect 15051 1516 15085 1550
rect 14840 1425 14874 1459
rect 14915 1414 14949 1448
rect 14983 1419 15017 1453
rect 15051 1443 15085 1477
rect 14840 1357 14874 1391
rect 14915 1341 14949 1375
rect 14983 1346 15017 1380
rect 15051 1370 15085 1404
rect 14840 1289 14874 1323
rect 14915 1268 14949 1302
rect 14983 1273 15017 1307
rect 15051 1297 15085 1331
rect 14840 1221 14874 1255
rect 14915 1195 14949 1229
rect 14983 1200 15017 1234
rect 15051 1224 15085 1258
rect 14840 1153 14874 1187
rect 14915 1122 14949 1156
rect 14983 1127 15017 1161
rect 15051 1151 15085 1185
rect 14840 1085 14874 1119
rect 14840 1017 14874 1051
rect 14915 1049 14949 1083
rect 14983 1054 15017 1088
rect 15051 1078 15085 1112
rect 14840 949 14874 983
rect 14915 976 14949 1010
rect 14983 981 15017 1015
rect 15051 1005 15085 1039
rect 14840 881 14874 915
rect 14915 903 14949 937
rect 14983 908 15017 942
rect 15051 932 15085 966
rect 14840 813 14874 847
rect 14915 830 14949 864
rect 14983 835 15017 869
rect 15051 859 15085 893
rect 14840 745 14874 779
rect 14915 757 14949 791
rect 14983 762 15017 796
rect 15051 786 15085 820
rect 14840 677 14874 711
rect 14915 684 14949 718
rect 14983 689 15017 723
rect 15051 713 15085 747
rect 51 576 85 610
rect 119 576 153 610
rect 187 576 221 610
rect 262 609 296 643
rect 262 541 296 575
rect 51 504 85 538
rect 119 504 153 538
rect 187 504 221 538
rect 14840 609 14874 643
rect 14915 611 14949 645
rect 14983 616 15017 650
rect 15051 640 15085 674
rect 14840 541 14874 575
rect 14915 538 14949 572
rect 14983 543 15017 577
rect 15051 567 15085 601
rect 51 432 85 466
rect 119 432 153 466
rect 187 432 221 466
rect 302 465 336 499
rect 375 465 409 499
rect 448 465 482 499
rect 521 465 555 499
rect 594 465 628 499
rect 667 465 701 499
rect 740 465 774 499
rect 813 465 847 499
rect 886 465 920 499
rect 959 465 993 499
rect 1032 465 1066 499
rect 1105 465 1139 499
rect 1178 465 1212 499
rect 1251 465 1285 499
rect 1324 465 1358 499
rect 1397 465 1431 499
rect 1470 465 1504 499
rect 1543 465 1577 499
rect 1616 465 1650 499
rect 1689 465 1723 499
rect 1762 465 1796 499
rect 1835 465 1869 499
rect 1908 465 1942 499
rect 1981 465 2015 499
rect 2054 465 2088 499
rect 2127 465 2161 499
rect 2200 465 2234 499
rect 2273 465 2307 499
rect 2346 465 2380 499
rect 2419 465 2453 499
rect 2492 465 2526 499
rect 2565 465 2599 499
rect 2638 465 2672 499
rect 2711 465 2745 499
rect 2784 465 2818 499
rect 2857 465 2891 499
rect 2930 465 2964 499
rect 3003 465 3037 499
rect 3076 465 3110 499
rect 3149 465 3183 499
rect 3222 465 3256 499
rect 3295 465 3329 499
rect 3368 465 3402 499
rect 3441 465 3475 499
rect 3514 465 3548 499
rect 3587 465 3621 499
rect 3660 465 3694 499
rect 3733 465 3767 499
rect 3806 465 3840 499
rect 3879 465 3913 499
rect 3952 465 3986 499
rect 4025 465 4059 499
rect 4098 465 4132 499
rect 4171 465 4205 499
rect 4244 465 4278 499
rect 4317 465 4351 499
rect 4390 465 4424 499
rect 4463 465 4497 499
rect 4536 465 4570 499
rect 4609 465 4643 499
rect 4682 465 4716 499
rect 4755 465 4789 499
rect 4828 465 4862 499
rect 4901 465 4935 499
rect 4974 465 5008 499
rect 5047 465 5081 499
rect 5120 465 5154 499
rect 5193 465 5227 499
rect 5266 465 5300 499
rect 5339 465 5373 499
rect 5411 465 5445 499
rect 5483 465 5517 499
rect 5555 465 5589 499
rect 5627 465 5661 499
rect 5699 465 5733 499
rect 5771 465 5805 499
rect 5843 465 5877 499
rect 5915 465 5949 499
rect 5987 465 6021 499
rect 6059 465 6093 499
rect 6131 465 6165 499
rect 6203 465 6237 499
rect 6275 465 6309 499
rect 6347 465 6381 499
rect 6419 465 6453 499
rect 6491 465 6525 499
rect 6563 465 6597 499
rect 6635 465 6669 499
rect 6707 465 6741 499
rect 6779 465 6813 499
rect 6851 465 6885 499
rect 6923 465 6957 499
rect 6995 465 7029 499
rect 7067 465 7101 499
rect 7139 465 7173 499
rect 7211 465 7245 499
rect 7283 465 7317 499
rect 7355 465 7389 499
rect 7427 465 7461 499
rect 7499 465 7533 499
rect 7571 465 7605 499
rect 7643 465 7677 499
rect 7715 465 7749 499
rect 7787 465 7821 499
rect 7859 465 7893 499
rect 7931 465 7965 499
rect 8003 465 8037 499
rect 8075 465 8109 499
rect 8147 465 8181 499
rect 8219 465 8253 499
rect 8291 465 8325 499
rect 8363 465 8397 499
rect 8435 465 8469 499
rect 8507 465 8541 499
rect 8579 465 8613 499
rect 8651 465 8685 499
rect 8723 465 8757 499
rect 8795 465 8829 499
rect 8867 465 8901 499
rect 8939 465 8973 499
rect 9011 465 9045 499
rect 9083 465 9117 499
rect 9155 465 9189 499
rect 9227 465 9261 499
rect 9299 465 9333 499
rect 9371 465 9405 499
rect 9443 465 9477 499
rect 9515 465 9549 499
rect 9587 465 9621 499
rect 9659 465 9693 499
rect 9731 465 9765 499
rect 9803 465 9837 499
rect 9875 465 9909 499
rect 9947 465 9981 499
rect 10019 465 10053 499
rect 10091 465 10125 499
rect 10163 465 10197 499
rect 10235 465 10269 499
rect 10307 465 10341 499
rect 10379 465 10413 499
rect 10451 465 10485 499
rect 10523 465 10557 499
rect 10595 465 10629 499
rect 10667 465 10701 499
rect 10739 465 10773 499
rect 10811 465 10845 499
rect 10883 465 10917 499
rect 10955 465 10989 499
rect 11027 465 11061 499
rect 11099 465 11133 499
rect 11171 465 11205 499
rect 11243 465 11277 499
rect 11315 465 11349 499
rect 11387 465 11421 499
rect 11459 465 11493 499
rect 11531 465 11565 499
rect 11603 465 11637 499
rect 11675 465 11709 499
rect 11747 465 11781 499
rect 11819 465 11853 499
rect 11891 465 11925 499
rect 11963 465 11997 499
rect 12035 465 12069 499
rect 12107 465 12141 499
rect 12179 465 12213 499
rect 12251 465 12285 499
rect 12323 465 12357 499
rect 12395 465 12429 499
rect 12467 465 12501 499
rect 12539 465 12573 499
rect 12611 465 12645 499
rect 12683 465 12717 499
rect 12755 465 12789 499
rect 12827 465 12861 499
rect 12899 465 12933 499
rect 12971 465 13005 499
rect 13043 465 13077 499
rect 13115 465 13149 499
rect 13187 465 13221 499
rect 13259 465 13293 499
rect 13331 465 13365 499
rect 13403 465 13437 499
rect 13475 465 13509 499
rect 13547 465 13581 499
rect 13619 465 13653 499
rect 13691 465 13725 499
rect 13763 465 13797 499
rect 13835 465 13869 499
rect 13907 465 13941 499
rect 13979 465 14013 499
rect 14051 465 14085 499
rect 14123 465 14157 499
rect 14195 465 14229 499
rect 14267 465 14301 499
rect 14339 465 14373 499
rect 14411 465 14445 499
rect 14483 465 14517 499
rect 14555 465 14589 499
rect 14627 465 14661 499
rect 14699 465 14733 499
rect 14771 465 14805 499
rect 14843 465 14877 499
rect 14915 465 14949 499
rect 14983 470 15017 504
rect 15051 494 15085 528
rect 302 397 336 431
rect 375 397 409 431
rect 448 397 482 431
rect 521 397 555 431
rect 594 397 628 431
rect 667 397 701 431
rect 740 397 774 431
rect 813 397 847 431
rect 886 397 920 431
rect 959 397 993 431
rect 1032 397 1066 431
rect 1105 397 1139 431
rect 1178 397 1212 431
rect 1251 397 1285 431
rect 1324 397 1358 431
rect 1397 397 1431 431
rect 1470 397 1504 431
rect 1543 397 1577 431
rect 1616 397 1650 431
rect 1689 397 1723 431
rect 1762 397 1796 431
rect 1835 397 1869 431
rect 1908 397 1942 431
rect 1981 397 2015 431
rect 2054 397 2088 431
rect 2127 397 2161 431
rect 2200 397 2234 431
rect 2273 397 2307 431
rect 2346 397 2380 431
rect 2419 397 2453 431
rect 2492 397 2526 431
rect 2565 397 2599 431
rect 2638 397 2672 431
rect 2711 397 2745 431
rect 2784 397 2818 431
rect 2857 397 2891 431
rect 2930 397 2964 431
rect 3003 397 3037 431
rect 3076 397 3110 431
rect 3149 397 3183 431
rect 3222 397 3256 431
rect 3295 397 3329 431
rect 3368 397 3402 431
rect 3441 397 3475 431
rect 3514 397 3548 431
rect 3587 397 3621 431
rect 3660 397 3694 431
rect 3733 397 3767 431
rect 3806 397 3840 431
rect 3879 397 3913 431
rect 3952 397 3986 431
rect 4025 397 4059 431
rect 4098 397 4132 431
rect 4171 397 4205 431
rect 4244 397 4278 431
rect 4317 397 4351 431
rect 4390 397 4424 431
rect 4463 397 4497 431
rect 4536 397 4570 431
rect 4609 397 4643 431
rect 4682 397 4716 431
rect 4755 397 4789 431
rect 4828 397 4862 431
rect 4901 397 4935 431
rect 4974 397 5008 431
rect 5047 397 5081 431
rect 5119 397 5153 431
rect 5191 397 5225 431
rect 5263 397 5297 431
rect 5335 397 5369 431
rect 5407 397 5441 431
rect 5479 397 5513 431
rect 5551 397 5585 431
rect 5623 397 5657 431
rect 5695 397 5729 431
rect 5767 397 5801 431
rect 5839 397 5873 431
rect 5911 397 5945 431
rect 5983 397 6017 431
rect 6055 397 6089 431
rect 6127 397 6161 431
rect 6199 397 6233 431
rect 6271 397 6305 431
rect 6343 397 6377 431
rect 6415 397 6449 431
rect 6487 397 6521 431
rect 6559 397 6593 431
rect 6631 397 6665 431
rect 6703 397 6737 431
rect 6775 397 6809 431
rect 6847 397 6881 431
rect 6919 397 6953 431
rect 6991 397 7025 431
rect 7063 397 7097 431
rect 7135 397 7169 431
rect 7207 397 7241 431
rect 7279 397 7313 431
rect 7351 397 7385 431
rect 7423 397 7457 431
rect 7495 397 7529 431
rect 7567 397 7601 431
rect 7639 397 7673 431
rect 7711 397 7745 431
rect 7783 397 7817 431
rect 7855 397 7889 431
rect 7927 397 7961 431
rect 7999 397 8033 431
rect 8071 397 8105 431
rect 8143 397 8177 431
rect 8215 397 8249 431
rect 8287 397 8321 431
rect 8359 397 8393 431
rect 8431 397 8465 431
rect 8503 397 8537 431
rect 8575 397 8609 431
rect 8647 397 8681 431
rect 8719 397 8753 431
rect 8791 397 8825 431
rect 8863 397 8897 431
rect 8935 397 8969 431
rect 9007 397 9041 431
rect 9079 397 9113 431
rect 9151 397 9185 431
rect 9223 397 9257 431
rect 9295 397 9329 431
rect 9367 397 9401 431
rect 9439 397 9473 431
rect 9511 397 9545 431
rect 9583 397 9617 431
rect 9655 397 9689 431
rect 9727 397 9761 431
rect 9799 397 9833 431
rect 9871 397 9905 431
rect 9943 397 9977 431
rect 10015 397 10049 431
rect 10087 397 10121 431
rect 10159 397 10193 431
rect 10231 397 10265 431
rect 10303 397 10337 431
rect 10375 397 10409 431
rect 10447 397 10481 431
rect 10519 397 10553 431
rect 10591 397 10625 431
rect 10663 397 10697 431
rect 10735 397 10769 431
rect 10807 397 10841 431
rect 10879 397 10913 431
rect 10951 397 10985 431
rect 11023 397 11057 431
rect 11095 397 11129 431
rect 11167 397 11201 431
rect 11239 397 11273 431
rect 11311 397 11345 431
rect 11383 397 11417 431
rect 11455 397 11489 431
rect 11527 397 11561 431
rect 11599 397 11633 431
rect 11671 397 11705 431
rect 11743 397 11777 431
rect 11815 397 11849 431
rect 11887 397 11921 431
rect 11959 397 11993 431
rect 12031 397 12065 431
rect 12103 397 12137 431
rect 12175 397 12209 431
rect 12247 397 12281 431
rect 12319 397 12353 431
rect 12391 397 12425 431
rect 12463 397 12497 431
rect 12535 397 12569 431
rect 12607 397 12641 431
rect 12679 397 12713 431
rect 12751 397 12785 431
rect 12823 397 12857 431
rect 12895 397 12929 431
rect 12967 397 13001 431
rect 13039 397 13073 431
rect 13111 397 13145 431
rect 13183 397 13217 431
rect 13255 397 13289 431
rect 13327 397 13361 431
rect 13399 397 13433 431
rect 13471 397 13505 431
rect 13543 397 13577 431
rect 13615 397 13649 431
rect 13687 397 13721 431
rect 13759 397 13793 431
rect 13831 397 13865 431
rect 13903 397 13937 431
rect 13975 397 14009 431
rect 14047 397 14081 431
rect 14119 397 14153 431
rect 14191 397 14225 431
rect 14263 397 14297 431
rect 14335 397 14369 431
rect 14407 397 14441 431
rect 14479 397 14513 431
rect 14551 397 14585 431
rect 14623 397 14657 431
rect 14695 397 14729 431
rect 14767 397 14801 431
rect 14839 397 14873 431
rect 14911 397 14945 431
rect 14983 397 15017 431
rect 15051 421 15085 455
rect 51 360 85 394
rect 119 360 153 394
rect 187 360 221 394
rect 302 329 336 363
rect 375 329 409 363
rect 448 329 482 363
rect 521 329 555 363
rect 594 329 628 363
rect 667 329 701 363
rect 740 329 774 363
rect 813 329 847 363
rect 886 329 920 363
rect 959 329 993 363
rect 1032 329 1066 363
rect 1105 329 1139 363
rect 1178 329 1212 363
rect 1251 329 1285 363
rect 1324 329 1358 363
rect 1397 329 1431 363
rect 1470 329 1504 363
rect 1543 329 1577 363
rect 1616 329 1650 363
rect 1689 329 1723 363
rect 1762 329 1796 363
rect 1835 329 1869 363
rect 1908 329 1942 363
rect 1981 329 2015 363
rect 2054 329 2088 363
rect 2127 329 2161 363
rect 2200 329 2234 363
rect 2273 329 2307 363
rect 2346 329 2380 363
rect 2419 329 2453 363
rect 2492 329 2526 363
rect 2565 329 2599 363
rect 2638 329 2672 363
rect 2711 329 2745 363
rect 2784 329 2818 363
rect 2857 329 2891 363
rect 2930 329 2964 363
rect 3003 329 3037 363
rect 3076 329 3110 363
rect 3149 329 3183 363
rect 3222 329 3256 363
rect 3295 329 3329 363
rect 3368 329 3402 363
rect 3440 329 3474 363
rect 3512 329 3546 363
rect 3584 329 3618 363
rect 3656 329 3690 363
rect 3728 329 3762 363
rect 3800 329 3834 363
rect 3872 329 3906 363
rect 3944 329 3978 363
rect 4016 329 4050 363
rect 4088 329 4122 363
rect 4160 329 4194 363
rect 4232 329 4266 363
rect 4304 329 4338 363
rect 4376 329 4410 363
rect 4448 329 4482 363
rect 4520 329 4554 363
rect 4592 329 4626 363
rect 4664 329 4698 363
rect 4736 329 4770 363
rect 4808 329 4842 363
rect 4880 329 4914 363
rect 4952 329 4986 363
rect 5024 329 5058 363
rect 5096 329 5130 363
rect 5168 329 5202 363
rect 5240 329 5274 363
rect 5312 329 5346 363
rect 5384 329 5418 363
rect 5456 329 5490 363
rect 5528 329 5562 363
rect 5600 329 5634 363
rect 5672 329 5706 363
rect 5744 329 5778 363
rect 5816 329 5850 363
rect 5888 329 5922 363
rect 5960 329 5994 363
rect 6032 329 6066 363
rect 6104 329 6138 363
rect 6176 329 6210 363
rect 6248 329 6282 363
rect 6320 329 6354 363
rect 6392 329 6426 363
rect 6464 329 6498 363
rect 6536 329 6570 363
rect 6608 329 6642 363
rect 6680 329 6714 363
rect 6752 329 6786 363
rect 6824 329 6858 363
rect 6896 329 6930 363
rect 6968 329 7002 363
rect 7040 329 7074 363
rect 7112 329 7146 363
rect 7184 329 7218 363
rect 7256 329 7290 363
rect 7328 329 7362 363
rect 7400 329 7434 363
rect 7472 329 7506 363
rect 7544 329 7578 363
rect 7616 329 7650 363
rect 7688 329 7722 363
rect 7760 329 7794 363
rect 7832 329 7866 363
rect 7904 329 7938 363
rect 7976 329 8010 363
rect 8048 329 8082 363
rect 8120 329 8154 363
rect 8192 329 8226 363
rect 8264 329 8298 363
rect 8336 329 8370 363
rect 8408 329 8442 363
rect 8480 329 8514 363
rect 8552 329 8586 363
rect 8624 329 8658 363
rect 8696 329 8730 363
rect 8768 329 8802 363
rect 8840 329 8874 363
rect 8912 329 8946 363
rect 8984 329 9018 363
rect 9056 329 9090 363
rect 9128 329 9162 363
rect 9200 329 9234 363
rect 9272 329 9306 363
rect 9344 329 9378 363
rect 9416 329 9450 363
rect 9488 329 9522 363
rect 9560 329 9594 363
rect 9632 329 9666 363
rect 9704 329 9738 363
rect 9776 329 9810 363
rect 9848 329 9882 363
rect 9920 329 9954 363
rect 9992 329 10026 363
rect 10064 329 10098 363
rect 10136 329 10170 363
rect 10208 329 10242 363
rect 10280 329 10314 363
rect 10352 329 10386 363
rect 10424 329 10458 363
rect 10496 329 10530 363
rect 10568 329 10602 363
rect 10640 329 10674 363
rect 10712 329 10746 363
rect 10784 329 10818 363
rect 10856 329 10890 363
rect 10928 329 10962 363
rect 11000 329 11034 363
rect 11072 329 11106 363
rect 11144 329 11178 363
rect 11216 329 11250 363
rect 11288 329 11322 363
rect 11360 329 11394 363
rect 11432 329 11466 363
rect 11504 329 11538 363
rect 11576 329 11610 363
rect 11648 329 11682 363
rect 11720 329 11754 363
rect 11792 329 11826 363
rect 11864 329 11898 363
rect 11936 329 11970 363
rect 12008 329 12042 363
rect 12080 329 12114 363
rect 12152 329 12186 363
rect 12224 329 12258 363
rect 12296 329 12330 363
rect 12368 329 12402 363
rect 12440 329 12474 363
rect 12512 329 12546 363
rect 12584 329 12618 363
rect 12656 329 12690 363
rect 12728 329 12762 363
rect 12800 329 12834 363
rect 12872 329 12906 363
rect 12944 329 12978 363
rect 13016 329 13050 363
rect 13088 329 13122 363
rect 13160 329 13194 363
rect 13232 329 13266 363
rect 13304 329 13338 363
rect 13376 329 13410 363
rect 13448 329 13482 363
rect 13520 329 13554 363
rect 13592 329 13626 363
rect 13664 329 13698 363
rect 13736 329 13770 363
rect 13808 329 13842 363
rect 13880 329 13914 363
rect 13952 329 13986 363
rect 14024 329 14058 363
rect 14096 329 14130 363
rect 14168 329 14202 363
rect 14240 329 14274 363
rect 14312 329 14346 363
rect 14384 329 14418 363
rect 14456 329 14490 363
rect 14528 329 14562 363
rect 14600 329 14634 363
rect 14672 329 14706 363
rect 14744 329 14778 363
rect 14816 329 14850 363
rect 14888 329 14922 363
rect 14960 329 14994 363
rect 15051 348 15085 382
<< mvnsubdiffcont >>
rect 497 4585 531 4619
rect 584 4570 10410 4638
rect 10445 4604 10479 4638
rect 10514 4604 10548 4638
rect 10583 4604 10617 4638
rect 10652 4604 10686 4638
rect 10721 4604 10755 4638
rect 10790 4604 10824 4638
rect 10859 4604 10893 4638
rect 10928 4604 10962 4638
rect 10997 4604 11031 4638
rect 11066 4604 11100 4638
rect 11135 4604 11169 4638
rect 11204 4604 11238 4638
rect 11273 4604 11307 4638
rect 11342 4604 11376 4638
rect 11411 4604 11445 4638
rect 11480 4604 11514 4638
rect 11549 4604 11583 4638
rect 11618 4604 11652 4638
rect 11687 4604 11721 4638
rect 11756 4604 11790 4638
rect 11825 4604 11859 4638
rect 11894 4604 11928 4638
rect 11963 4604 11997 4638
rect 12032 4604 12066 4638
rect 12101 4604 12135 4638
rect 12170 4604 12204 4638
rect 12239 4604 12273 4638
rect 12308 4604 12342 4638
rect 12377 4604 12411 4638
rect 12446 4604 12480 4638
rect 12515 4604 12549 4638
rect 12584 4604 12618 4638
rect 12653 4604 12687 4638
rect 12722 4604 12756 4638
rect 12791 4604 12825 4638
rect 12860 4604 12894 4638
rect 12929 4604 12963 4638
rect 12998 4604 13032 4638
rect 13067 4604 13101 4638
rect 13136 4604 13170 4638
rect 13205 4604 13239 4638
rect 13274 4604 13308 4638
rect 13343 4604 13377 4638
rect 13412 4604 13446 4638
rect 13481 4604 13515 4638
rect 13550 4604 13584 4638
rect 13619 4604 13653 4638
rect 13688 4604 13722 4638
rect 13757 4604 13791 4638
rect 13826 4604 13860 4638
rect 13895 4604 13929 4638
rect 13964 4604 13998 4638
rect 14033 4604 14067 4638
rect 14102 4604 14136 4638
rect 14171 4604 14205 4638
rect 14240 4604 14274 4638
rect 14309 4604 14343 4638
rect 14378 4604 14412 4638
rect 14447 4604 14481 4638
rect 14516 4604 14550 4638
rect 14585 4604 14619 4638
rect 497 4515 531 4549
rect 565 4536 12363 4570
rect 12397 4536 12431 4570
rect 12466 4536 12500 4570
rect 12535 4536 12569 4570
rect 12604 4536 12638 4570
rect 12673 4536 12707 4570
rect 12742 4536 12776 4570
rect 12811 4536 12845 4570
rect 12880 4536 12914 4570
rect 12949 4536 12983 4570
rect 13018 4536 13052 4570
rect 13087 4536 13121 4570
rect 13156 4536 13190 4570
rect 13225 4536 13259 4570
rect 13294 4536 13328 4570
rect 13363 4536 13397 4570
rect 13432 4536 13466 4570
rect 13501 4536 13535 4570
rect 13570 4536 13604 4570
rect 13639 4536 13673 4570
rect 13708 4536 13742 4570
rect 13777 4536 13811 4570
rect 13846 4536 13880 4570
rect 13915 4536 13949 4570
rect 13984 4536 14018 4570
rect 14053 4536 14087 4570
rect 14122 4536 14156 4570
rect 14191 4536 14225 4570
rect 14260 4536 14294 4570
rect 14329 4536 14363 4570
rect 14398 4536 14432 4570
rect 14467 4536 14501 4570
rect 14536 4551 14570 4570
rect 497 4445 531 4479
rect 565 4464 599 4498
rect 633 4468 12363 4536
rect 14536 4502 14638 4551
rect 12398 4468 12432 4502
rect 12467 4468 12501 4502
rect 12536 4468 12570 4502
rect 12605 4468 12639 4502
rect 12674 4468 12708 4502
rect 12743 4468 12777 4502
rect 12812 4468 12846 4502
rect 12881 4468 12915 4502
rect 12950 4468 12984 4502
rect 13019 4468 13053 4502
rect 13088 4468 13122 4502
rect 13157 4468 13191 4502
rect 13226 4468 13260 4502
rect 13295 4468 13329 4502
rect 13364 4468 13398 4502
rect 13433 4468 13467 4502
rect 13502 4468 13536 4502
rect 13571 4468 13605 4502
rect 13640 4468 13674 4502
rect 13709 4468 13743 4502
rect 13778 4468 13812 4502
rect 13847 4468 13881 4502
rect 13916 4468 13950 4502
rect 13985 4468 14019 4502
rect 14054 4468 14088 4502
rect 14123 4468 14157 4502
rect 14192 4468 14226 4502
rect 14261 4468 14295 4502
rect 14330 4468 14364 4502
rect 14399 4468 14433 4502
rect 497 4375 531 4409
rect 565 4392 599 4426
rect 633 4395 667 4429
rect 497 4305 531 4339
rect 565 4320 599 4354
rect 633 4322 667 4356
rect 497 4235 531 4269
rect 565 4248 599 4282
rect 633 4249 667 4283
rect 497 4165 531 4199
rect 565 4176 599 4210
rect 633 4177 667 4211
rect 497 4095 531 4129
rect 565 4104 599 4138
rect 633 4105 667 4139
rect 497 4025 531 4059
rect 565 4032 599 4066
rect 633 4033 667 4067
rect 497 3955 531 3989
rect 565 3960 599 3994
rect 633 3961 667 3995
rect 497 3886 531 3920
rect 565 3888 599 3922
rect 633 3889 667 3923
rect 497 3817 531 3851
rect 565 3817 599 3851
rect 633 3817 667 3851
rect 497 3715 531 3749
rect 565 3715 599 3749
rect 633 3715 667 3749
rect 497 3646 531 3680
rect 565 3646 599 3680
rect 633 3646 667 3680
rect 497 3577 531 3611
rect 565 3577 599 3611
rect 633 3577 667 3611
rect 497 3508 531 3542
rect 565 3508 599 3542
rect 633 3508 667 3542
rect 497 3439 531 3473
rect 565 3439 599 3473
rect 633 3439 667 3473
rect 497 3370 531 3404
rect 565 3370 599 3404
rect 633 3370 667 3404
rect 497 3301 531 3335
rect 565 3301 599 3335
rect 633 3301 667 3335
rect 497 3232 531 3266
rect 565 3232 599 3266
rect 633 3232 667 3266
rect 497 3163 531 3197
rect 565 3163 599 3197
rect 633 3163 667 3197
rect 1635 4048 1669 4082
rect 1635 3980 1669 4014
rect 1635 3912 1669 3946
rect 1635 3844 1669 3878
rect 1635 3776 1669 3810
rect 1635 3708 1669 3742
rect 1635 3640 1669 3674
rect 1635 3572 1669 3606
rect 1635 3504 1669 3538
rect 1635 3436 1669 3470
rect 1635 3368 1669 3402
rect 1635 3300 1669 3334
rect 1635 3232 1669 3266
rect 1635 3164 1669 3198
rect 2627 4048 2661 4082
rect 2627 3980 2661 4014
rect 2627 3912 2661 3946
rect 2627 3844 2661 3878
rect 2627 3776 2661 3810
rect 2627 3708 2661 3742
rect 2627 3640 2661 3674
rect 2627 3572 2661 3606
rect 2627 3504 2661 3538
rect 2627 3436 2661 3470
rect 2627 3368 2661 3402
rect 2627 3300 2661 3334
rect 2627 3232 2661 3266
rect 2627 3164 2661 3198
rect 3619 4048 3653 4082
rect 3619 3980 3653 4014
rect 3619 3912 3653 3946
rect 3619 3844 3653 3878
rect 3619 3776 3653 3810
rect 3619 3708 3653 3742
rect 3619 3640 3653 3674
rect 3619 3572 3653 3606
rect 3619 3504 3653 3538
rect 3619 3436 3653 3470
rect 3619 3368 3653 3402
rect 3619 3300 3653 3334
rect 3619 3232 3653 3266
rect 3619 3164 3653 3198
rect 4611 4048 4645 4082
rect 4611 3980 4645 4014
rect 4611 3912 4645 3946
rect 4611 3844 4645 3878
rect 4611 3776 4645 3810
rect 4611 3708 4645 3742
rect 4611 3640 4645 3674
rect 4611 3572 4645 3606
rect 4611 3504 4645 3538
rect 4611 3436 4645 3470
rect 4611 3368 4645 3402
rect 4611 3300 4645 3334
rect 4611 3232 4645 3266
rect 4611 3164 4645 3198
rect 5603 4048 5637 4082
rect 5603 3980 5637 4014
rect 5603 3912 5637 3946
rect 5603 3844 5637 3878
rect 5603 3776 5637 3810
rect 5603 3708 5637 3742
rect 5603 3640 5637 3674
rect 5603 3572 5637 3606
rect 5603 3504 5637 3538
rect 5603 3436 5637 3470
rect 5603 3368 5637 3402
rect 5603 3300 5637 3334
rect 5603 3232 5637 3266
rect 5603 3164 5637 3198
rect 6595 4048 6629 4082
rect 6595 3980 6629 4014
rect 6595 3912 6629 3946
rect 6595 3844 6629 3878
rect 6595 3776 6629 3810
rect 6595 3708 6629 3742
rect 6595 3640 6629 3674
rect 6595 3572 6629 3606
rect 6595 3504 6629 3538
rect 6595 3436 6629 3470
rect 6595 3368 6629 3402
rect 6595 3300 6629 3334
rect 6595 3232 6629 3266
rect 6595 3164 6629 3198
rect 7587 4048 7621 4082
rect 7587 3980 7621 4014
rect 7587 3912 7621 3946
rect 7587 3844 7621 3878
rect 7587 3776 7621 3810
rect 7587 3708 7621 3742
rect 7587 3640 7621 3674
rect 7587 3572 7621 3606
rect 7587 3504 7621 3538
rect 7587 3436 7621 3470
rect 7587 3368 7621 3402
rect 7587 3300 7621 3334
rect 7587 3232 7621 3266
rect 7587 3164 7621 3198
rect 8579 4048 8613 4082
rect 8579 3980 8613 4014
rect 8579 3912 8613 3946
rect 8579 3844 8613 3878
rect 8579 3776 8613 3810
rect 8579 3708 8613 3742
rect 8579 3640 8613 3674
rect 8579 3572 8613 3606
rect 8579 3504 8613 3538
rect 8579 3436 8613 3470
rect 8579 3368 8613 3402
rect 8579 3300 8613 3334
rect 8579 3232 8613 3266
rect 8579 3164 8613 3198
rect 9571 4048 9605 4082
rect 9571 3980 9605 4014
rect 9571 3912 9605 3946
rect 9571 3844 9605 3878
rect 9571 3776 9605 3810
rect 9571 3708 9605 3742
rect 9571 3640 9605 3674
rect 9571 3572 9605 3606
rect 9571 3504 9605 3538
rect 9571 3436 9605 3470
rect 9571 3368 9605 3402
rect 9571 3300 9605 3334
rect 9571 3232 9605 3266
rect 9571 3164 9605 3198
rect 10563 4048 10597 4082
rect 10563 3980 10597 4014
rect 10563 3912 10597 3946
rect 10563 3844 10597 3878
rect 10563 3776 10597 3810
rect 10563 3708 10597 3742
rect 10563 3640 10597 3674
rect 10563 3572 10597 3606
rect 10563 3504 10597 3538
rect 10563 3436 10597 3470
rect 10563 3368 10597 3402
rect 10563 3300 10597 3334
rect 10563 3232 10597 3266
rect 10563 3164 10597 3198
rect 11555 4048 11589 4082
rect 11555 3980 11589 4014
rect 11555 3912 11589 3946
rect 11555 3844 11589 3878
rect 11555 3776 11589 3810
rect 11555 3708 11589 3742
rect 11555 3640 11589 3674
rect 11555 3572 11589 3606
rect 11555 3504 11589 3538
rect 11555 3436 11589 3470
rect 11555 3368 11589 3402
rect 11555 3300 11589 3334
rect 11555 3232 11589 3266
rect 11555 3164 11589 3198
rect 12547 4048 12581 4082
rect 12547 3980 12581 4014
rect 12547 3912 12581 3946
rect 12547 3844 12581 3878
rect 12547 3776 12581 3810
rect 12547 3708 12581 3742
rect 12547 3640 12581 3674
rect 12547 3572 12581 3606
rect 12547 3504 12581 3538
rect 12547 3436 12581 3470
rect 12547 3368 12581 3402
rect 12547 3300 12581 3334
rect 12547 3232 12581 3266
rect 12547 3164 12581 3198
rect 13539 4048 13573 4082
rect 13539 3980 13573 4014
rect 13539 3912 13573 3946
rect 13539 3844 13573 3878
rect 13539 3776 13573 3810
rect 13539 3708 13573 3742
rect 13539 3640 13573 3674
rect 13539 3572 13573 3606
rect 13539 3504 13573 3538
rect 13539 3436 13573 3470
rect 13539 3368 13573 3402
rect 13539 3300 13573 3334
rect 13539 3232 13573 3266
rect 13539 3164 13573 3198
rect 14468 3992 14638 4502
rect 14468 3923 14502 3957
rect 14536 3924 14638 3992
rect 14604 3905 14638 3924
rect 14468 3854 14502 3888
rect 14536 3855 14570 3889
rect 14604 3837 14638 3871
rect 14468 3785 14502 3819
rect 14536 3786 14570 3820
rect 14604 3769 14638 3803
rect 14468 3716 14502 3750
rect 14536 3717 14570 3751
rect 14604 3701 14638 3735
rect 14468 3647 14502 3681
rect 14536 3648 14570 3682
rect 14604 3633 14638 3667
rect 14468 3578 14502 3612
rect 14536 3579 14570 3613
rect 14604 3565 14638 3599
rect 14468 3509 14502 3543
rect 14536 3510 14570 3544
rect 14604 3497 14638 3531
rect 14468 3440 14502 3474
rect 14536 3441 14570 3475
rect 14604 3429 14638 3463
rect 14468 3371 14502 3405
rect 14536 3372 14570 3406
rect 14604 3361 14638 3395
rect 14468 3302 14502 3336
rect 14536 3303 14570 3337
rect 14604 3293 14638 3327
rect 14468 3233 14502 3267
rect 14536 3234 14570 3268
rect 14604 3225 14638 3259
rect 14468 3164 14502 3198
rect 14536 3165 14570 3199
rect 14604 3157 14638 3191
rect 497 3094 531 3128
rect 565 3094 599 3128
rect 633 3094 667 3128
rect 497 3025 531 3059
rect 565 3025 599 3059
rect 633 3025 667 3059
rect 497 2956 531 2990
rect 565 2956 599 2990
rect 633 2956 667 2990
rect 497 2887 531 2921
rect 565 2887 599 2921
rect 633 2887 667 2921
rect 497 2818 531 2852
rect 565 2818 599 2852
rect 633 2818 667 2852
rect 497 2749 531 2783
rect 565 2749 599 2783
rect 633 2749 667 2783
rect 497 2680 531 2714
rect 565 2680 599 2714
rect 633 2680 667 2714
rect 497 2611 531 2645
rect 565 2611 599 2645
rect 633 2611 667 2645
rect 497 2542 531 2576
rect 565 2542 599 2576
rect 633 2542 667 2576
rect 1601 3010 1635 3044
rect 1669 3010 1703 3044
rect 1601 2940 1635 2974
rect 1669 2940 1703 2974
rect 1601 2870 1635 2904
rect 1669 2870 1703 2904
rect 1601 2800 1635 2834
rect 1669 2800 1703 2834
rect 1601 2730 1635 2764
rect 1669 2730 1703 2764
rect 1601 2660 1635 2694
rect 1669 2660 1703 2694
rect 2593 3010 2627 3044
rect 2661 3010 2695 3044
rect 2593 2940 2627 2974
rect 2661 2940 2695 2974
rect 2593 2870 2627 2904
rect 2661 2870 2695 2904
rect 2593 2800 2627 2834
rect 2661 2800 2695 2834
rect 2593 2730 2627 2764
rect 2661 2730 2695 2764
rect 2593 2660 2627 2694
rect 2661 2660 2695 2694
rect 3585 3010 3619 3044
rect 3653 3010 3687 3044
rect 3585 2940 3619 2974
rect 3653 2940 3687 2974
rect 3585 2870 3619 2904
rect 3653 2870 3687 2904
rect 3585 2800 3619 2834
rect 3653 2800 3687 2834
rect 3585 2730 3619 2764
rect 3653 2730 3687 2764
rect 3585 2660 3619 2694
rect 3653 2660 3687 2694
rect 4577 3010 4611 3044
rect 4645 3010 4679 3044
rect 4577 2940 4611 2974
rect 4645 2940 4679 2974
rect 4577 2870 4611 2904
rect 4645 2870 4679 2904
rect 4577 2800 4611 2834
rect 4645 2800 4679 2834
rect 4577 2730 4611 2764
rect 4645 2730 4679 2764
rect 4577 2660 4611 2694
rect 4645 2660 4679 2694
rect 5569 3010 5603 3044
rect 5637 3010 5671 3044
rect 5569 2940 5603 2974
rect 5637 2940 5671 2974
rect 5569 2870 5603 2904
rect 5637 2870 5671 2904
rect 5569 2800 5603 2834
rect 5637 2800 5671 2834
rect 5569 2730 5603 2764
rect 5637 2730 5671 2764
rect 5569 2660 5603 2694
rect 5637 2660 5671 2694
rect 6561 3010 6595 3044
rect 6629 3010 6663 3044
rect 6561 2940 6595 2974
rect 6629 2940 6663 2974
rect 6561 2870 6595 2904
rect 6629 2870 6663 2904
rect 6561 2800 6595 2834
rect 6629 2800 6663 2834
rect 6561 2730 6595 2764
rect 6629 2730 6663 2764
rect 6561 2660 6595 2694
rect 6629 2660 6663 2694
rect 7553 3010 7587 3044
rect 7621 3010 7655 3044
rect 7553 2940 7587 2974
rect 7621 2940 7655 2974
rect 7553 2870 7587 2904
rect 7621 2870 7655 2904
rect 7553 2800 7587 2834
rect 7621 2800 7655 2834
rect 7553 2730 7587 2764
rect 7621 2730 7655 2764
rect 7553 2660 7587 2694
rect 7621 2660 7655 2694
rect 8545 3010 8579 3044
rect 8613 3010 8647 3044
rect 8545 2940 8579 2974
rect 8613 2940 8647 2974
rect 8545 2870 8579 2904
rect 8613 2870 8647 2904
rect 8545 2800 8579 2834
rect 8613 2800 8647 2834
rect 8545 2730 8579 2764
rect 8613 2730 8647 2764
rect 8545 2660 8579 2694
rect 8613 2660 8647 2694
rect 9537 3010 9571 3044
rect 9605 3010 9639 3044
rect 9537 2940 9571 2974
rect 9605 2940 9639 2974
rect 9537 2870 9571 2904
rect 9605 2870 9639 2904
rect 9537 2800 9571 2834
rect 9605 2800 9639 2834
rect 9537 2730 9571 2764
rect 9605 2730 9639 2764
rect 9537 2660 9571 2694
rect 9605 2660 9639 2694
rect 10529 3010 10563 3044
rect 10597 3010 10631 3044
rect 10529 2940 10563 2974
rect 10597 2940 10631 2974
rect 10529 2870 10563 2904
rect 10597 2870 10631 2904
rect 10529 2800 10563 2834
rect 10597 2800 10631 2834
rect 10529 2730 10563 2764
rect 10597 2730 10631 2764
rect 10529 2660 10563 2694
rect 10597 2660 10631 2694
rect 11521 3010 11555 3044
rect 11589 3010 11623 3044
rect 11521 2940 11555 2974
rect 11589 2940 11623 2974
rect 11521 2870 11555 2904
rect 11589 2870 11623 2904
rect 11521 2800 11555 2834
rect 11589 2800 11623 2834
rect 11521 2730 11555 2764
rect 11589 2730 11623 2764
rect 11521 2660 11555 2694
rect 11589 2660 11623 2694
rect 12513 3010 12547 3044
rect 12581 3010 12615 3044
rect 12513 2940 12547 2974
rect 12581 2940 12615 2974
rect 12513 2870 12547 2904
rect 12581 2870 12615 2904
rect 12513 2800 12547 2834
rect 12581 2800 12615 2834
rect 12513 2730 12547 2764
rect 12581 2730 12615 2764
rect 12513 2660 12547 2694
rect 12581 2660 12615 2694
rect 13505 3010 13539 3044
rect 13573 3010 13607 3044
rect 13505 2940 13539 2974
rect 13573 2940 13607 2974
rect 13505 2870 13539 2904
rect 13573 2870 13607 2904
rect 13505 2800 13539 2834
rect 13573 2800 13607 2834
rect 13505 2730 13539 2764
rect 13573 2730 13607 2764
rect 13505 2660 13539 2694
rect 13573 2660 13607 2694
rect 14468 3095 14502 3129
rect 14536 3096 14570 3130
rect 14604 3089 14638 3123
rect 14468 3026 14502 3060
rect 14536 3027 14570 3061
rect 14604 3021 14638 3055
rect 14468 2957 14502 2991
rect 14536 2958 14570 2992
rect 14604 2953 14638 2987
rect 14468 2888 14502 2922
rect 14536 2889 14570 2923
rect 14604 2885 14638 2919
rect 14468 2819 14502 2853
rect 14536 2820 14570 2854
rect 14604 2817 14638 2851
rect 14468 2750 14502 2784
rect 14536 2751 14570 2785
rect 14604 2749 14638 2783
rect 14468 2681 14502 2715
rect 14536 2682 14570 2716
rect 14604 2681 14638 2715
rect 14468 2612 14502 2646
rect 14536 2613 14570 2647
rect 14604 2613 14638 2647
rect 497 2473 531 2507
rect 565 2473 599 2507
rect 633 2473 667 2507
rect 497 2404 531 2438
rect 565 2404 599 2438
rect 633 2404 667 2438
rect 497 2335 531 2369
rect 565 2335 599 2369
rect 633 2335 667 2369
rect 497 2266 531 2300
rect 565 2266 599 2300
rect 633 2266 667 2300
rect 497 2197 531 2231
rect 565 2197 599 2231
rect 633 2197 667 2231
rect 497 2129 531 2163
rect 565 2128 599 2162
rect 633 2128 667 2162
rect 497 2061 531 2095
rect 565 2059 599 2093
rect 633 2059 667 2093
rect 497 1993 531 2027
rect 565 1990 599 2024
rect 633 1990 667 2024
rect 497 1925 531 1959
rect 565 1921 599 1955
rect 633 1921 667 1955
rect 497 1857 531 1891
rect 565 1852 599 1886
rect 633 1852 667 1886
rect 497 1789 531 1823
rect 565 1783 599 1817
rect 633 1783 667 1817
rect 497 1721 531 1755
rect 565 1714 599 1748
rect 633 1714 667 1748
rect 497 1653 531 1687
rect 565 1645 599 1679
rect 633 1645 667 1679
rect 497 1585 531 1619
rect 565 1576 599 1610
rect 633 1576 667 1610
rect 1635 2506 1669 2540
rect 1635 2438 1669 2472
rect 1635 2370 1669 2404
rect 1635 2302 1669 2336
rect 1635 2234 1669 2268
rect 1635 2166 1669 2200
rect 1635 2098 1669 2132
rect 1635 2030 1669 2064
rect 1635 1962 1669 1996
rect 1635 1894 1669 1928
rect 1635 1826 1669 1860
rect 1635 1758 1669 1792
rect 1635 1690 1669 1724
rect 1635 1622 1669 1656
rect 2627 2506 2661 2540
rect 2627 2438 2661 2472
rect 2627 2370 2661 2404
rect 2627 2302 2661 2336
rect 2627 2234 2661 2268
rect 2627 2166 2661 2200
rect 2627 2098 2661 2132
rect 2627 2030 2661 2064
rect 2627 1962 2661 1996
rect 2627 1894 2661 1928
rect 2627 1826 2661 1860
rect 2627 1758 2661 1792
rect 2627 1690 2661 1724
rect 2627 1622 2661 1656
rect 3619 2506 3653 2540
rect 3619 2438 3653 2472
rect 3619 2370 3653 2404
rect 3619 2302 3653 2336
rect 3619 2234 3653 2268
rect 3619 2166 3653 2200
rect 3619 2098 3653 2132
rect 3619 2030 3653 2064
rect 3619 1962 3653 1996
rect 3619 1894 3653 1928
rect 3619 1826 3653 1860
rect 3619 1758 3653 1792
rect 3619 1690 3653 1724
rect 3619 1622 3653 1656
rect 4611 2506 4645 2540
rect 4611 2438 4645 2472
rect 4611 2370 4645 2404
rect 4611 2302 4645 2336
rect 4611 2234 4645 2268
rect 4611 2166 4645 2200
rect 4611 2098 4645 2132
rect 4611 2030 4645 2064
rect 4611 1962 4645 1996
rect 4611 1894 4645 1928
rect 4611 1826 4645 1860
rect 4611 1758 4645 1792
rect 4611 1690 4645 1724
rect 4611 1622 4645 1656
rect 5603 2506 5637 2540
rect 5603 2438 5637 2472
rect 5603 2370 5637 2404
rect 5603 2302 5637 2336
rect 5603 2234 5637 2268
rect 5603 2166 5637 2200
rect 5603 2098 5637 2132
rect 5603 2030 5637 2064
rect 5603 1962 5637 1996
rect 5603 1894 5637 1928
rect 5603 1826 5637 1860
rect 5603 1758 5637 1792
rect 5603 1690 5637 1724
rect 5603 1622 5637 1656
rect 6595 2506 6629 2540
rect 6595 2438 6629 2472
rect 6595 2370 6629 2404
rect 6595 2302 6629 2336
rect 6595 2234 6629 2268
rect 6595 2166 6629 2200
rect 6595 2098 6629 2132
rect 6595 2030 6629 2064
rect 6595 1962 6629 1996
rect 6595 1894 6629 1928
rect 6595 1826 6629 1860
rect 6595 1758 6629 1792
rect 6595 1690 6629 1724
rect 6595 1622 6629 1656
rect 7587 2506 7621 2540
rect 7587 2438 7621 2472
rect 7587 2370 7621 2404
rect 7587 2302 7621 2336
rect 7587 2234 7621 2268
rect 7587 2166 7621 2200
rect 7587 2098 7621 2132
rect 7587 2030 7621 2064
rect 7587 1962 7621 1996
rect 7587 1894 7621 1928
rect 7587 1826 7621 1860
rect 7587 1758 7621 1792
rect 7587 1690 7621 1724
rect 7587 1622 7621 1656
rect 8579 2506 8613 2540
rect 8579 2438 8613 2472
rect 8579 2370 8613 2404
rect 8579 2302 8613 2336
rect 8579 2234 8613 2268
rect 8579 2166 8613 2200
rect 8579 2098 8613 2132
rect 8579 2030 8613 2064
rect 8579 1962 8613 1996
rect 8579 1894 8613 1928
rect 8579 1826 8613 1860
rect 8579 1758 8613 1792
rect 8579 1690 8613 1724
rect 8579 1622 8613 1656
rect 9571 2506 9605 2540
rect 9571 2438 9605 2472
rect 9571 2370 9605 2404
rect 9571 2302 9605 2336
rect 9571 2234 9605 2268
rect 9571 2166 9605 2200
rect 9571 2098 9605 2132
rect 9571 2030 9605 2064
rect 9571 1962 9605 1996
rect 9571 1894 9605 1928
rect 9571 1826 9605 1860
rect 9571 1758 9605 1792
rect 9571 1690 9605 1724
rect 9571 1622 9605 1656
rect 10563 2506 10597 2540
rect 10563 2438 10597 2472
rect 10563 2370 10597 2404
rect 10563 2302 10597 2336
rect 10563 2234 10597 2268
rect 10563 2166 10597 2200
rect 10563 2098 10597 2132
rect 10563 2030 10597 2064
rect 10563 1962 10597 1996
rect 10563 1894 10597 1928
rect 10563 1826 10597 1860
rect 10563 1758 10597 1792
rect 10563 1690 10597 1724
rect 10563 1622 10597 1656
rect 11555 2506 11589 2540
rect 11555 2438 11589 2472
rect 11555 2370 11589 2404
rect 11555 2302 11589 2336
rect 11555 2234 11589 2268
rect 11555 2166 11589 2200
rect 11555 2098 11589 2132
rect 11555 2030 11589 2064
rect 11555 1962 11589 1996
rect 11555 1894 11589 1928
rect 11555 1826 11589 1860
rect 11555 1758 11589 1792
rect 11555 1690 11589 1724
rect 11555 1622 11589 1656
rect 12547 2506 12581 2540
rect 12547 2438 12581 2472
rect 12547 2370 12581 2404
rect 12547 2302 12581 2336
rect 12547 2234 12581 2268
rect 12547 2166 12581 2200
rect 12547 2098 12581 2132
rect 12547 2030 12581 2064
rect 12547 1962 12581 1996
rect 12547 1894 12581 1928
rect 12547 1826 12581 1860
rect 12547 1758 12581 1792
rect 12547 1690 12581 1724
rect 12547 1622 12581 1656
rect 13539 2506 13573 2540
rect 13539 2438 13573 2472
rect 13539 2370 13573 2404
rect 13539 2302 13573 2336
rect 13539 2234 13573 2268
rect 13539 2166 13573 2200
rect 13539 2098 13573 2132
rect 13539 2030 13573 2064
rect 13539 1962 13573 1996
rect 13539 1894 13573 1928
rect 13539 1826 13573 1860
rect 13539 1758 13573 1792
rect 13539 1690 13573 1724
rect 13539 1622 13573 1656
rect 14468 2543 14502 2577
rect 14536 2544 14570 2578
rect 14604 2545 14638 2579
rect 14468 2474 14502 2508
rect 14536 2475 14570 2509
rect 14604 2477 14638 2511
rect 14468 2405 14502 2439
rect 14536 2406 14570 2440
rect 14604 2409 14638 2443
rect 14468 2336 14502 2370
rect 14536 2337 14570 2371
rect 14604 2341 14638 2375
rect 14468 2267 14502 2301
rect 14536 2268 14570 2302
rect 14604 2273 14638 2307
rect 14468 2198 14502 2232
rect 14536 2199 14570 2233
rect 14604 2205 14638 2239
rect 14468 2129 14502 2163
rect 14536 2130 14570 2164
rect 14604 2137 14638 2171
rect 14468 2060 14502 2094
rect 14536 2061 14570 2095
rect 14604 2069 14638 2103
rect 14468 1991 14502 2025
rect 14536 1992 14570 2026
rect 14604 2001 14638 2035
rect 14468 1922 14502 1956
rect 14536 1923 14570 1957
rect 14604 1933 14638 1967
rect 14468 1853 14502 1887
rect 14536 1854 14570 1888
rect 14604 1865 14638 1899
rect 14468 1784 14502 1818
rect 14536 1785 14570 1819
rect 14604 1797 14638 1831
rect 14468 1715 14502 1749
rect 14536 1716 14570 1750
rect 14604 1729 14638 1763
rect 14468 1646 14502 1680
rect 14536 1647 14570 1681
rect 14604 1661 14638 1695
rect 14468 1577 14502 1611
rect 14536 1578 14570 1612
rect 14604 1593 14638 1627
rect 497 1517 531 1551
rect 565 1507 599 1541
rect 633 1507 667 1541
rect 497 1449 531 1483
rect 565 1438 599 1472
rect 633 1438 667 1472
rect 497 1381 531 1415
rect 565 1369 599 1403
rect 633 1369 667 1403
rect 14468 1508 14502 1542
rect 14536 1509 14570 1543
rect 14604 1525 14638 1559
rect 14468 1439 14502 1473
rect 14536 1440 14570 1474
rect 14604 1457 14638 1491
rect 497 1313 531 1347
rect 565 1300 599 1334
rect 633 1300 667 1334
rect 497 1245 531 1279
rect 565 1231 599 1265
rect 633 1231 667 1265
rect 497 1177 531 1211
rect 565 1162 599 1196
rect 633 1162 667 1196
rect 497 1109 531 1143
rect 565 1093 599 1127
rect 633 1093 667 1127
rect 497 1041 531 1075
rect 565 1024 599 1058
rect 633 1024 667 1058
rect 497 973 531 1007
rect 565 955 599 989
rect 633 955 667 989
rect 497 920 531 939
rect 497 818 667 920
rect 14468 1370 14502 1404
rect 14536 1371 14570 1405
rect 14604 1389 14638 1423
rect 14468 1301 14502 1335
rect 14536 1302 14570 1336
rect 14604 1321 14638 1355
rect 14468 1232 14502 1266
rect 14536 1233 14570 1267
rect 14604 1253 14638 1287
rect 14468 1163 14502 1197
rect 14536 1164 14570 1198
rect 14604 1184 14638 1218
rect 14468 1094 14502 1128
rect 14536 1095 14570 1129
rect 14604 1115 14638 1149
rect 14468 1025 14502 1059
rect 14536 1026 14570 1060
rect 14604 1046 14638 1080
rect 14468 956 14502 990
rect 14536 957 14570 991
rect 14604 977 14638 1011
rect 14468 887 14502 921
rect 14536 888 14570 922
rect 14604 908 14638 942
rect 702 818 736 852
rect 771 818 805 852
rect 840 818 874 852
rect 909 818 943 852
rect 978 818 1012 852
rect 1047 818 1081 852
rect 1116 818 1150 852
rect 1185 818 1219 852
rect 1254 818 1288 852
rect 1323 818 1357 852
rect 1392 818 1426 852
rect 1461 818 1495 852
rect 1530 818 1564 852
rect 1599 818 1633 852
rect 1668 818 1702 852
rect 1737 818 1771 852
rect 1806 818 1840 852
rect 1875 818 1909 852
rect 1944 818 1978 852
rect 2013 818 2047 852
rect 2082 818 2116 852
rect 2151 818 2185 852
rect 2220 818 2254 852
rect 2289 818 2323 852
rect 2358 818 2392 852
rect 2427 818 2461 852
rect 2496 818 2530 852
rect 2565 818 2599 852
rect 2634 818 2668 852
rect 2703 818 2737 852
rect 497 769 599 818
rect 2772 784 14502 852
rect 14536 819 14570 853
rect 14604 839 14638 873
rect 565 750 599 769
rect 634 750 668 784
rect 703 750 737 784
rect 772 750 806 784
rect 841 750 875 784
rect 910 750 944 784
rect 979 750 1013 784
rect 1048 750 1082 784
rect 1117 750 1151 784
rect 1186 750 1220 784
rect 1255 750 1289 784
rect 1324 750 1358 784
rect 1393 750 1427 784
rect 1462 750 1496 784
rect 1531 750 1565 784
rect 1600 750 1634 784
rect 1669 750 1703 784
rect 1738 750 1772 784
rect 1807 750 1841 784
rect 1876 750 1910 784
rect 1945 750 1979 784
rect 2014 750 2048 784
rect 2083 750 2117 784
rect 2152 750 2186 784
rect 2221 750 2255 784
rect 2290 750 2324 784
rect 2359 750 2393 784
rect 2428 750 2462 784
rect 2497 750 2531 784
rect 2566 750 2600 784
rect 2635 750 2669 784
rect 2704 750 2738 784
rect 2772 750 14570 784
rect 14604 770 14638 804
rect 516 682 550 716
rect 585 682 619 716
rect 654 682 688 716
rect 723 682 757 716
rect 792 682 826 716
rect 861 682 895 716
rect 930 682 964 716
rect 999 682 1033 716
rect 1068 682 1102 716
rect 1137 682 1171 716
rect 1206 682 1240 716
rect 1275 682 1309 716
rect 1344 682 1378 716
rect 1413 682 1447 716
rect 1482 682 1516 716
rect 1551 682 1585 716
rect 1620 682 1654 716
rect 1689 682 1723 716
rect 1758 682 1792 716
rect 1827 682 1861 716
rect 1896 682 1930 716
rect 1965 682 1999 716
rect 2034 682 2068 716
rect 2103 682 2137 716
rect 2172 682 2206 716
rect 2241 682 2275 716
rect 2310 682 2344 716
rect 2379 682 2413 716
rect 2448 682 2482 716
rect 2517 682 2551 716
rect 2586 682 2620 716
rect 2655 682 2689 716
rect 2724 682 2758 716
rect 2793 682 2827 716
rect 2862 682 2896 716
rect 2931 682 2965 716
rect 3000 682 3034 716
rect 3069 682 3103 716
rect 3138 682 3172 716
rect 3207 682 3241 716
rect 3276 682 3310 716
rect 3345 682 3379 716
rect 3414 682 3448 716
rect 3483 682 3517 716
rect 3552 682 3586 716
rect 3621 682 3655 716
rect 3690 682 3724 716
rect 3759 682 3793 716
rect 3828 682 3862 716
rect 3897 682 3931 716
rect 3966 682 4000 716
rect 4035 682 4069 716
rect 4104 682 4138 716
rect 4173 682 4207 716
rect 4242 682 4276 716
rect 4311 682 4345 716
rect 4380 682 4414 716
rect 4449 682 4483 716
rect 4518 682 4552 716
rect 4587 682 4621 716
rect 4656 682 4690 716
rect 4725 682 14551 750
rect 14604 701 14638 735
<< poly >>
rect 881 4308 1001 4324
rect 881 4274 924 4308
rect 958 4274 1001 4308
rect 881 4234 1001 4274
rect 881 4200 924 4234
rect 958 4200 1001 4234
rect 881 4152 1001 4200
rect 1311 4308 1431 4324
rect 1311 4274 1354 4308
rect 1388 4274 1431 4308
rect 1311 4234 1431 4274
rect 1311 4200 1354 4234
rect 1388 4200 1431 4234
rect 1311 4152 1431 4200
rect 1873 4308 1993 4324
rect 1873 4274 1916 4308
rect 1950 4274 1993 4308
rect 1873 4234 1993 4274
rect 1873 4200 1916 4234
rect 1950 4200 1993 4234
rect 1873 4152 1993 4200
rect 2303 4308 2423 4324
rect 2303 4274 2346 4308
rect 2380 4274 2423 4308
rect 2303 4234 2423 4274
rect 2303 4200 2346 4234
rect 2380 4200 2423 4234
rect 2303 4152 2423 4200
rect 2865 4308 2985 4324
rect 2865 4274 2908 4308
rect 2942 4274 2985 4308
rect 2865 4234 2985 4274
rect 2865 4200 2908 4234
rect 2942 4200 2985 4234
rect 2865 4152 2985 4200
rect 3295 4308 3415 4324
rect 3295 4274 3338 4308
rect 3372 4274 3415 4308
rect 3295 4234 3415 4274
rect 3295 4200 3338 4234
rect 3372 4200 3415 4234
rect 3295 4152 3415 4200
rect 3857 4308 3977 4324
rect 3857 4274 3900 4308
rect 3934 4274 3977 4308
rect 3857 4234 3977 4274
rect 3857 4200 3900 4234
rect 3934 4200 3977 4234
rect 3857 4152 3977 4200
rect 4287 4308 4407 4324
rect 4287 4274 4330 4308
rect 4364 4274 4407 4308
rect 4287 4234 4407 4274
rect 4287 4200 4330 4234
rect 4364 4200 4407 4234
rect 4287 4152 4407 4200
rect 4849 4308 4969 4324
rect 4849 4274 4892 4308
rect 4926 4274 4969 4308
rect 4849 4234 4969 4274
rect 4849 4200 4892 4234
rect 4926 4200 4969 4234
rect 4849 4152 4969 4200
rect 5279 4308 5399 4324
rect 5279 4274 5322 4308
rect 5356 4274 5399 4308
rect 5279 4234 5399 4274
rect 5279 4200 5322 4234
rect 5356 4200 5399 4234
rect 5279 4152 5399 4200
rect 5841 4308 5961 4324
rect 5841 4274 5884 4308
rect 5918 4274 5961 4308
rect 5841 4234 5961 4274
rect 5841 4200 5884 4234
rect 5918 4200 5961 4234
rect 5841 4152 5961 4200
rect 6271 4308 6391 4324
rect 6271 4274 6314 4308
rect 6348 4274 6391 4308
rect 6271 4234 6391 4274
rect 6271 4200 6314 4234
rect 6348 4200 6391 4234
rect 6271 4152 6391 4200
rect 6833 4308 6953 4324
rect 6833 4274 6876 4308
rect 6910 4274 6953 4308
rect 6833 4234 6953 4274
rect 6833 4200 6876 4234
rect 6910 4200 6953 4234
rect 6833 4152 6953 4200
rect 7263 4308 7383 4324
rect 7263 4274 7306 4308
rect 7340 4274 7383 4308
rect 7263 4234 7383 4274
rect 7263 4200 7306 4234
rect 7340 4200 7383 4234
rect 7263 4152 7383 4200
rect 7825 4308 7945 4324
rect 7825 4274 7868 4308
rect 7902 4274 7945 4308
rect 7825 4234 7945 4274
rect 7825 4200 7868 4234
rect 7902 4200 7945 4234
rect 7825 4152 7945 4200
rect 8255 4308 8375 4324
rect 8255 4274 8298 4308
rect 8332 4274 8375 4308
rect 8255 4234 8375 4274
rect 8255 4200 8298 4234
rect 8332 4200 8375 4234
rect 8255 4152 8375 4200
rect 8817 4308 8937 4324
rect 8817 4274 8860 4308
rect 8894 4274 8937 4308
rect 8817 4234 8937 4274
rect 8817 4200 8860 4234
rect 8894 4200 8937 4234
rect 8817 4152 8937 4200
rect 9247 4308 9367 4324
rect 9247 4274 9290 4308
rect 9324 4274 9367 4308
rect 9247 4234 9367 4274
rect 9247 4200 9290 4234
rect 9324 4200 9367 4234
rect 9247 4152 9367 4200
rect 9809 4308 9929 4324
rect 9809 4274 9852 4308
rect 9886 4274 9929 4308
rect 9809 4234 9929 4274
rect 9809 4200 9852 4234
rect 9886 4200 9929 4234
rect 9809 4152 9929 4200
rect 10239 4308 10359 4324
rect 10239 4274 10282 4308
rect 10316 4274 10359 4308
rect 10239 4234 10359 4274
rect 10239 4200 10282 4234
rect 10316 4200 10359 4234
rect 10239 4152 10359 4200
rect 10801 4308 10921 4324
rect 10801 4274 10844 4308
rect 10878 4274 10921 4308
rect 10801 4234 10921 4274
rect 10801 4200 10844 4234
rect 10878 4200 10921 4234
rect 10801 4152 10921 4200
rect 11231 4308 11351 4324
rect 11231 4274 11274 4308
rect 11308 4274 11351 4308
rect 11231 4234 11351 4274
rect 11231 4200 11274 4234
rect 11308 4200 11351 4234
rect 11231 4152 11351 4200
rect 11793 4308 11913 4324
rect 11793 4274 11836 4308
rect 11870 4274 11913 4308
rect 11793 4234 11913 4274
rect 11793 4200 11836 4234
rect 11870 4200 11913 4234
rect 11793 4152 11913 4200
rect 12223 4308 12343 4324
rect 12223 4274 12266 4308
rect 12300 4274 12343 4308
rect 12223 4234 12343 4274
rect 12223 4200 12266 4234
rect 12300 4200 12343 4234
rect 12223 4152 12343 4200
rect 12785 4308 12905 4324
rect 12785 4274 12828 4308
rect 12862 4274 12905 4308
rect 12785 4234 12905 4274
rect 12785 4200 12828 4234
rect 12862 4200 12905 4234
rect 12785 4152 12905 4200
rect 13215 4308 13335 4324
rect 13215 4274 13258 4308
rect 13292 4274 13335 4308
rect 13215 4234 13335 4274
rect 13215 4200 13258 4234
rect 13292 4200 13335 4234
rect 13215 4152 13335 4200
rect 13777 4308 13897 4324
rect 13777 4274 13820 4308
rect 13854 4274 13897 4308
rect 13777 4234 13897 4274
rect 13777 4200 13820 4234
rect 13854 4200 13897 4234
rect 13777 4152 13897 4200
rect 14135 4308 14255 4324
rect 14135 4274 14178 4308
rect 14212 4274 14255 4308
rect 14135 4234 14255 4274
rect 14135 4200 14178 4234
rect 14212 4200 14255 4234
rect 14135 4152 14255 4200
rect 881 3104 1001 3152
rect 881 3070 924 3104
rect 958 3070 1001 3104
rect 881 3026 1001 3070
rect 881 2992 924 3026
rect 958 2992 1001 3026
rect 881 2948 1001 2992
rect 881 2914 924 2948
rect 958 2914 1001 2948
rect 881 2870 1001 2914
rect 881 2836 924 2870
rect 958 2836 1001 2870
rect 881 2792 1001 2836
rect 881 2758 924 2792
rect 958 2758 1001 2792
rect 881 2713 1001 2758
rect 881 2679 924 2713
rect 958 2679 1001 2713
rect 881 2634 1001 2679
rect 881 2600 924 2634
rect 958 2600 1001 2634
rect 881 2552 1001 2600
rect 1311 3104 1431 3152
rect 1311 3070 1354 3104
rect 1388 3070 1431 3104
rect 1873 3104 1993 3152
rect 1311 3026 1431 3070
rect 1311 2992 1354 3026
rect 1388 2992 1431 3026
rect 1311 2948 1431 2992
rect 1311 2914 1354 2948
rect 1388 2914 1431 2948
rect 1311 2870 1431 2914
rect 1311 2836 1354 2870
rect 1388 2836 1431 2870
rect 1311 2792 1431 2836
rect 1311 2758 1354 2792
rect 1388 2758 1431 2792
rect 1311 2713 1431 2758
rect 1311 2679 1354 2713
rect 1388 2679 1431 2713
rect 1311 2634 1431 2679
rect 1311 2600 1354 2634
rect 1388 2600 1431 2634
rect 1873 3070 1916 3104
rect 1950 3070 1993 3104
rect 1873 3026 1993 3070
rect 1873 2992 1916 3026
rect 1950 2992 1993 3026
rect 1873 2948 1993 2992
rect 1873 2914 1916 2948
rect 1950 2914 1993 2948
rect 1873 2870 1993 2914
rect 1873 2836 1916 2870
rect 1950 2836 1993 2870
rect 1873 2792 1993 2836
rect 1873 2758 1916 2792
rect 1950 2758 1993 2792
rect 1873 2713 1993 2758
rect 1873 2679 1916 2713
rect 1950 2679 1993 2713
rect 1873 2634 1993 2679
rect 1311 2552 1431 2600
rect 1873 2600 1916 2634
rect 1950 2600 1993 2634
rect 1873 2552 1993 2600
rect 2303 3104 2423 3152
rect 2303 3070 2346 3104
rect 2380 3070 2423 3104
rect 2865 3104 2985 3152
rect 2303 3026 2423 3070
rect 2303 2992 2346 3026
rect 2380 2992 2423 3026
rect 2303 2948 2423 2992
rect 2303 2914 2346 2948
rect 2380 2914 2423 2948
rect 2303 2870 2423 2914
rect 2303 2836 2346 2870
rect 2380 2836 2423 2870
rect 2303 2792 2423 2836
rect 2303 2758 2346 2792
rect 2380 2758 2423 2792
rect 2303 2713 2423 2758
rect 2303 2679 2346 2713
rect 2380 2679 2423 2713
rect 2303 2634 2423 2679
rect 2303 2600 2346 2634
rect 2380 2600 2423 2634
rect 2865 3070 2908 3104
rect 2942 3070 2985 3104
rect 2865 3026 2985 3070
rect 2865 2992 2908 3026
rect 2942 2992 2985 3026
rect 2865 2948 2985 2992
rect 2865 2914 2908 2948
rect 2942 2914 2985 2948
rect 2865 2870 2985 2914
rect 2865 2836 2908 2870
rect 2942 2836 2985 2870
rect 2865 2792 2985 2836
rect 2865 2758 2908 2792
rect 2942 2758 2985 2792
rect 2865 2713 2985 2758
rect 2865 2679 2908 2713
rect 2942 2679 2985 2713
rect 2865 2634 2985 2679
rect 2303 2552 2423 2600
rect 2865 2600 2908 2634
rect 2942 2600 2985 2634
rect 2865 2552 2985 2600
rect 3295 3104 3415 3152
rect 3295 3070 3338 3104
rect 3372 3070 3415 3104
rect 3857 3104 3977 3152
rect 3295 3026 3415 3070
rect 3295 2992 3338 3026
rect 3372 2992 3415 3026
rect 3295 2948 3415 2992
rect 3295 2914 3338 2948
rect 3372 2914 3415 2948
rect 3295 2870 3415 2914
rect 3295 2836 3338 2870
rect 3372 2836 3415 2870
rect 3295 2792 3415 2836
rect 3295 2758 3338 2792
rect 3372 2758 3415 2792
rect 3295 2713 3415 2758
rect 3295 2679 3338 2713
rect 3372 2679 3415 2713
rect 3295 2634 3415 2679
rect 3295 2600 3338 2634
rect 3372 2600 3415 2634
rect 3857 3070 3900 3104
rect 3934 3070 3977 3104
rect 3857 3026 3977 3070
rect 3857 2992 3900 3026
rect 3934 2992 3977 3026
rect 3857 2948 3977 2992
rect 3857 2914 3900 2948
rect 3934 2914 3977 2948
rect 3857 2870 3977 2914
rect 3857 2836 3900 2870
rect 3934 2836 3977 2870
rect 3857 2792 3977 2836
rect 3857 2758 3900 2792
rect 3934 2758 3977 2792
rect 3857 2713 3977 2758
rect 3857 2679 3900 2713
rect 3934 2679 3977 2713
rect 3857 2634 3977 2679
rect 3295 2552 3415 2600
rect 3857 2600 3900 2634
rect 3934 2600 3977 2634
rect 3857 2552 3977 2600
rect 4287 3104 4407 3152
rect 4287 3070 4330 3104
rect 4364 3070 4407 3104
rect 4849 3104 4969 3152
rect 4287 3026 4407 3070
rect 4287 2992 4330 3026
rect 4364 2992 4407 3026
rect 4287 2948 4407 2992
rect 4287 2914 4330 2948
rect 4364 2914 4407 2948
rect 4287 2870 4407 2914
rect 4287 2836 4330 2870
rect 4364 2836 4407 2870
rect 4287 2792 4407 2836
rect 4287 2758 4330 2792
rect 4364 2758 4407 2792
rect 4287 2713 4407 2758
rect 4287 2679 4330 2713
rect 4364 2679 4407 2713
rect 4287 2634 4407 2679
rect 4287 2600 4330 2634
rect 4364 2600 4407 2634
rect 4849 3070 4892 3104
rect 4926 3070 4969 3104
rect 4849 3026 4969 3070
rect 4849 2992 4892 3026
rect 4926 2992 4969 3026
rect 4849 2948 4969 2992
rect 4849 2914 4892 2948
rect 4926 2914 4969 2948
rect 4849 2870 4969 2914
rect 4849 2836 4892 2870
rect 4926 2836 4969 2870
rect 4849 2792 4969 2836
rect 4849 2758 4892 2792
rect 4926 2758 4969 2792
rect 4849 2713 4969 2758
rect 4849 2679 4892 2713
rect 4926 2679 4969 2713
rect 4849 2634 4969 2679
rect 4287 2552 4407 2600
rect 4849 2600 4892 2634
rect 4926 2600 4969 2634
rect 4849 2552 4969 2600
rect 5279 3104 5399 3152
rect 5279 3070 5322 3104
rect 5356 3070 5399 3104
rect 5841 3104 5961 3152
rect 5279 3026 5399 3070
rect 5279 2992 5322 3026
rect 5356 2992 5399 3026
rect 5279 2948 5399 2992
rect 5279 2914 5322 2948
rect 5356 2914 5399 2948
rect 5279 2870 5399 2914
rect 5279 2836 5322 2870
rect 5356 2836 5399 2870
rect 5279 2792 5399 2836
rect 5279 2758 5322 2792
rect 5356 2758 5399 2792
rect 5279 2713 5399 2758
rect 5279 2679 5322 2713
rect 5356 2679 5399 2713
rect 5279 2634 5399 2679
rect 5279 2600 5322 2634
rect 5356 2600 5399 2634
rect 5841 3070 5884 3104
rect 5918 3070 5961 3104
rect 5841 3026 5961 3070
rect 5841 2992 5884 3026
rect 5918 2992 5961 3026
rect 5841 2948 5961 2992
rect 5841 2914 5884 2948
rect 5918 2914 5961 2948
rect 5841 2870 5961 2914
rect 5841 2836 5884 2870
rect 5918 2836 5961 2870
rect 5841 2792 5961 2836
rect 5841 2758 5884 2792
rect 5918 2758 5961 2792
rect 5841 2713 5961 2758
rect 5841 2679 5884 2713
rect 5918 2679 5961 2713
rect 5841 2634 5961 2679
rect 5279 2552 5399 2600
rect 5841 2600 5884 2634
rect 5918 2600 5961 2634
rect 5841 2552 5961 2600
rect 6271 3104 6391 3152
rect 6271 3070 6314 3104
rect 6348 3070 6391 3104
rect 6833 3104 6953 3152
rect 6271 3026 6391 3070
rect 6271 2992 6314 3026
rect 6348 2992 6391 3026
rect 6271 2948 6391 2992
rect 6271 2914 6314 2948
rect 6348 2914 6391 2948
rect 6271 2870 6391 2914
rect 6271 2836 6314 2870
rect 6348 2836 6391 2870
rect 6271 2792 6391 2836
rect 6271 2758 6314 2792
rect 6348 2758 6391 2792
rect 6271 2713 6391 2758
rect 6271 2679 6314 2713
rect 6348 2679 6391 2713
rect 6271 2634 6391 2679
rect 6271 2600 6314 2634
rect 6348 2600 6391 2634
rect 6833 3070 6876 3104
rect 6910 3070 6953 3104
rect 6833 3026 6953 3070
rect 6833 2992 6876 3026
rect 6910 2992 6953 3026
rect 6833 2948 6953 2992
rect 6833 2914 6876 2948
rect 6910 2914 6953 2948
rect 6833 2870 6953 2914
rect 6833 2836 6876 2870
rect 6910 2836 6953 2870
rect 6833 2792 6953 2836
rect 6833 2758 6876 2792
rect 6910 2758 6953 2792
rect 6833 2713 6953 2758
rect 6833 2679 6876 2713
rect 6910 2679 6953 2713
rect 6833 2634 6953 2679
rect 6271 2552 6391 2600
rect 6833 2600 6876 2634
rect 6910 2600 6953 2634
rect 6833 2552 6953 2600
rect 7263 3104 7383 3152
rect 7263 3070 7306 3104
rect 7340 3070 7383 3104
rect 7825 3104 7945 3152
rect 7263 3026 7383 3070
rect 7263 2992 7306 3026
rect 7340 2992 7383 3026
rect 7263 2948 7383 2992
rect 7263 2914 7306 2948
rect 7340 2914 7383 2948
rect 7263 2870 7383 2914
rect 7263 2836 7306 2870
rect 7340 2836 7383 2870
rect 7263 2792 7383 2836
rect 7263 2758 7306 2792
rect 7340 2758 7383 2792
rect 7263 2713 7383 2758
rect 7263 2679 7306 2713
rect 7340 2679 7383 2713
rect 7263 2634 7383 2679
rect 7263 2600 7306 2634
rect 7340 2600 7383 2634
rect 7825 3070 7868 3104
rect 7902 3070 7945 3104
rect 7825 3026 7945 3070
rect 7825 2992 7868 3026
rect 7902 2992 7945 3026
rect 7825 2948 7945 2992
rect 7825 2914 7868 2948
rect 7902 2914 7945 2948
rect 7825 2870 7945 2914
rect 7825 2836 7868 2870
rect 7902 2836 7945 2870
rect 7825 2792 7945 2836
rect 7825 2758 7868 2792
rect 7902 2758 7945 2792
rect 7825 2713 7945 2758
rect 7825 2679 7868 2713
rect 7902 2679 7945 2713
rect 7825 2634 7945 2679
rect 7263 2552 7383 2600
rect 7825 2600 7868 2634
rect 7902 2600 7945 2634
rect 7825 2552 7945 2600
rect 8255 3104 8375 3152
rect 8255 3070 8298 3104
rect 8332 3070 8375 3104
rect 8817 3104 8937 3152
rect 8255 3026 8375 3070
rect 8255 2992 8298 3026
rect 8332 2992 8375 3026
rect 8255 2948 8375 2992
rect 8255 2914 8298 2948
rect 8332 2914 8375 2948
rect 8255 2870 8375 2914
rect 8255 2836 8298 2870
rect 8332 2836 8375 2870
rect 8255 2792 8375 2836
rect 8255 2758 8298 2792
rect 8332 2758 8375 2792
rect 8255 2713 8375 2758
rect 8255 2679 8298 2713
rect 8332 2679 8375 2713
rect 8255 2634 8375 2679
rect 8255 2600 8298 2634
rect 8332 2600 8375 2634
rect 8817 3070 8860 3104
rect 8894 3070 8937 3104
rect 8817 3026 8937 3070
rect 8817 2992 8860 3026
rect 8894 2992 8937 3026
rect 8817 2948 8937 2992
rect 8817 2914 8860 2948
rect 8894 2914 8937 2948
rect 8817 2870 8937 2914
rect 8817 2836 8860 2870
rect 8894 2836 8937 2870
rect 8817 2792 8937 2836
rect 8817 2758 8860 2792
rect 8894 2758 8937 2792
rect 8817 2713 8937 2758
rect 8817 2679 8860 2713
rect 8894 2679 8937 2713
rect 8817 2634 8937 2679
rect 8255 2552 8375 2600
rect 8817 2600 8860 2634
rect 8894 2600 8937 2634
rect 8817 2552 8937 2600
rect 9247 3104 9367 3152
rect 9247 3070 9290 3104
rect 9324 3070 9367 3104
rect 9809 3104 9929 3152
rect 9247 3026 9367 3070
rect 9247 2992 9290 3026
rect 9324 2992 9367 3026
rect 9247 2948 9367 2992
rect 9247 2914 9290 2948
rect 9324 2914 9367 2948
rect 9247 2870 9367 2914
rect 9247 2836 9290 2870
rect 9324 2836 9367 2870
rect 9247 2792 9367 2836
rect 9247 2758 9290 2792
rect 9324 2758 9367 2792
rect 9247 2713 9367 2758
rect 9247 2679 9290 2713
rect 9324 2679 9367 2713
rect 9247 2634 9367 2679
rect 9247 2600 9290 2634
rect 9324 2600 9367 2634
rect 9809 3070 9852 3104
rect 9886 3070 9929 3104
rect 9809 3026 9929 3070
rect 9809 2992 9852 3026
rect 9886 2992 9929 3026
rect 9809 2948 9929 2992
rect 9809 2914 9852 2948
rect 9886 2914 9929 2948
rect 9809 2870 9929 2914
rect 9809 2836 9852 2870
rect 9886 2836 9929 2870
rect 9809 2792 9929 2836
rect 9809 2758 9852 2792
rect 9886 2758 9929 2792
rect 9809 2713 9929 2758
rect 9809 2679 9852 2713
rect 9886 2679 9929 2713
rect 9809 2634 9929 2679
rect 9247 2552 9367 2600
rect 9809 2600 9852 2634
rect 9886 2600 9929 2634
rect 9809 2552 9929 2600
rect 10239 3104 10359 3152
rect 10239 3070 10282 3104
rect 10316 3070 10359 3104
rect 10801 3104 10921 3152
rect 10239 3026 10359 3070
rect 10239 2992 10282 3026
rect 10316 2992 10359 3026
rect 10239 2948 10359 2992
rect 10239 2914 10282 2948
rect 10316 2914 10359 2948
rect 10239 2870 10359 2914
rect 10239 2836 10282 2870
rect 10316 2836 10359 2870
rect 10239 2792 10359 2836
rect 10239 2758 10282 2792
rect 10316 2758 10359 2792
rect 10239 2713 10359 2758
rect 10239 2679 10282 2713
rect 10316 2679 10359 2713
rect 10239 2634 10359 2679
rect 10239 2600 10282 2634
rect 10316 2600 10359 2634
rect 10801 3070 10844 3104
rect 10878 3070 10921 3104
rect 10801 3026 10921 3070
rect 10801 2992 10844 3026
rect 10878 2992 10921 3026
rect 10801 2948 10921 2992
rect 10801 2914 10844 2948
rect 10878 2914 10921 2948
rect 10801 2870 10921 2914
rect 10801 2836 10844 2870
rect 10878 2836 10921 2870
rect 10801 2792 10921 2836
rect 10801 2758 10844 2792
rect 10878 2758 10921 2792
rect 10801 2713 10921 2758
rect 10801 2679 10844 2713
rect 10878 2679 10921 2713
rect 10801 2634 10921 2679
rect 10239 2552 10359 2600
rect 10801 2600 10844 2634
rect 10878 2600 10921 2634
rect 10801 2552 10921 2600
rect 11231 3104 11351 3152
rect 11231 3070 11274 3104
rect 11308 3070 11351 3104
rect 11793 3104 11913 3152
rect 11231 3026 11351 3070
rect 11231 2992 11274 3026
rect 11308 2992 11351 3026
rect 11231 2948 11351 2992
rect 11231 2914 11274 2948
rect 11308 2914 11351 2948
rect 11231 2870 11351 2914
rect 11231 2836 11274 2870
rect 11308 2836 11351 2870
rect 11231 2792 11351 2836
rect 11231 2758 11274 2792
rect 11308 2758 11351 2792
rect 11231 2713 11351 2758
rect 11231 2679 11274 2713
rect 11308 2679 11351 2713
rect 11231 2634 11351 2679
rect 11231 2600 11274 2634
rect 11308 2600 11351 2634
rect 11793 3070 11836 3104
rect 11870 3070 11913 3104
rect 11793 3026 11913 3070
rect 11793 2992 11836 3026
rect 11870 2992 11913 3026
rect 11793 2948 11913 2992
rect 11793 2914 11836 2948
rect 11870 2914 11913 2948
rect 11793 2870 11913 2914
rect 11793 2836 11836 2870
rect 11870 2836 11913 2870
rect 11793 2792 11913 2836
rect 11793 2758 11836 2792
rect 11870 2758 11913 2792
rect 11793 2713 11913 2758
rect 11793 2679 11836 2713
rect 11870 2679 11913 2713
rect 11793 2634 11913 2679
rect 11231 2552 11351 2600
rect 11793 2600 11836 2634
rect 11870 2600 11913 2634
rect 11793 2552 11913 2600
rect 12223 3104 12343 3152
rect 12223 3070 12266 3104
rect 12300 3070 12343 3104
rect 12785 3104 12905 3152
rect 12223 3026 12343 3070
rect 12223 2992 12266 3026
rect 12300 2992 12343 3026
rect 12223 2948 12343 2992
rect 12223 2914 12266 2948
rect 12300 2914 12343 2948
rect 12223 2870 12343 2914
rect 12223 2836 12266 2870
rect 12300 2836 12343 2870
rect 12223 2792 12343 2836
rect 12223 2758 12266 2792
rect 12300 2758 12343 2792
rect 12223 2713 12343 2758
rect 12223 2679 12266 2713
rect 12300 2679 12343 2713
rect 12223 2634 12343 2679
rect 12223 2600 12266 2634
rect 12300 2600 12343 2634
rect 12785 3070 12828 3104
rect 12862 3070 12905 3104
rect 12785 3026 12905 3070
rect 12785 2992 12828 3026
rect 12862 2992 12905 3026
rect 12785 2948 12905 2992
rect 12785 2914 12828 2948
rect 12862 2914 12905 2948
rect 12785 2870 12905 2914
rect 12785 2836 12828 2870
rect 12862 2836 12905 2870
rect 12785 2792 12905 2836
rect 12785 2758 12828 2792
rect 12862 2758 12905 2792
rect 12785 2713 12905 2758
rect 12785 2679 12828 2713
rect 12862 2679 12905 2713
rect 12785 2634 12905 2679
rect 12223 2552 12343 2600
rect 12785 2600 12828 2634
rect 12862 2600 12905 2634
rect 12785 2552 12905 2600
rect 13215 3104 13335 3152
rect 13215 3070 13258 3104
rect 13292 3070 13335 3104
rect 13777 3104 13897 3152
rect 13215 3026 13335 3070
rect 13215 2992 13258 3026
rect 13292 2992 13335 3026
rect 13215 2948 13335 2992
rect 13215 2914 13258 2948
rect 13292 2914 13335 2948
rect 13215 2870 13335 2914
rect 13215 2836 13258 2870
rect 13292 2836 13335 2870
rect 13215 2792 13335 2836
rect 13215 2758 13258 2792
rect 13292 2758 13335 2792
rect 13215 2713 13335 2758
rect 13215 2679 13258 2713
rect 13292 2679 13335 2713
rect 13215 2634 13335 2679
rect 13215 2600 13258 2634
rect 13292 2600 13335 2634
rect 13777 3070 13820 3104
rect 13854 3070 13897 3104
rect 13777 3026 13897 3070
rect 13777 2992 13820 3026
rect 13854 2992 13897 3026
rect 13777 2948 13897 2992
rect 13777 2914 13820 2948
rect 13854 2914 13897 2948
rect 13777 2870 13897 2914
rect 13777 2836 13820 2870
rect 13854 2836 13897 2870
rect 13777 2792 13897 2836
rect 13777 2758 13820 2792
rect 13854 2758 13897 2792
rect 13777 2713 13897 2758
rect 13777 2679 13820 2713
rect 13854 2679 13897 2713
rect 13777 2634 13897 2679
rect 13215 2552 13335 2600
rect 13777 2600 13820 2634
rect 13854 2600 13897 2634
rect 13777 2552 13897 2600
rect 14135 3104 14255 3152
rect 14135 3070 14178 3104
rect 14212 3070 14255 3104
rect 14135 3026 14255 3070
rect 14135 2992 14178 3026
rect 14212 2992 14255 3026
rect 14135 2948 14255 2992
rect 14135 2914 14178 2948
rect 14212 2914 14255 2948
rect 14135 2870 14255 2914
rect 14135 2836 14178 2870
rect 14212 2836 14255 2870
rect 14135 2792 14255 2836
rect 14135 2758 14178 2792
rect 14212 2758 14255 2792
rect 14135 2713 14255 2758
rect 14135 2679 14178 2713
rect 14212 2679 14255 2713
rect 14135 2634 14255 2679
rect 14135 2600 14178 2634
rect 14212 2600 14255 2634
rect 14135 2552 14255 2600
rect 881 1504 1001 1552
rect 881 1470 924 1504
rect 958 1470 1001 1504
rect 881 1430 1001 1470
rect 881 1396 924 1430
rect 958 1396 1001 1430
rect 881 1380 1001 1396
rect 1311 1504 1431 1552
rect 1311 1470 1354 1504
rect 1388 1470 1431 1504
rect 1311 1430 1431 1470
rect 1311 1396 1354 1430
rect 1388 1396 1431 1430
rect 1311 1380 1431 1396
rect 1873 1504 1993 1552
rect 1873 1470 1916 1504
rect 1950 1470 1993 1504
rect 1873 1430 1993 1470
rect 1873 1396 1916 1430
rect 1950 1396 1993 1430
rect 1873 1380 1993 1396
rect 2303 1504 2423 1552
rect 2303 1470 2346 1504
rect 2380 1470 2423 1504
rect 2303 1430 2423 1470
rect 2303 1396 2346 1430
rect 2380 1396 2423 1430
rect 2303 1380 2423 1396
rect 2865 1504 2985 1552
rect 2865 1470 2908 1504
rect 2942 1470 2985 1504
rect 2865 1430 2985 1470
rect 2865 1396 2908 1430
rect 2942 1396 2985 1430
rect 2865 1380 2985 1396
rect 3295 1504 3415 1552
rect 3295 1470 3338 1504
rect 3372 1470 3415 1504
rect 3295 1430 3415 1470
rect 3295 1396 3338 1430
rect 3372 1396 3415 1430
rect 3295 1380 3415 1396
rect 3857 1504 3977 1552
rect 3857 1470 3900 1504
rect 3934 1470 3977 1504
rect 3857 1430 3977 1470
rect 3857 1396 3900 1430
rect 3934 1396 3977 1430
rect 3857 1380 3977 1396
rect 4287 1504 4407 1552
rect 4287 1470 4330 1504
rect 4364 1470 4407 1504
rect 4287 1430 4407 1470
rect 4287 1396 4330 1430
rect 4364 1396 4407 1430
rect 4287 1380 4407 1396
rect 4849 1504 4969 1552
rect 4849 1470 4892 1504
rect 4926 1470 4969 1504
rect 4849 1430 4969 1470
rect 4849 1396 4892 1430
rect 4926 1396 4969 1430
rect 4849 1380 4969 1396
rect 5279 1504 5399 1552
rect 5279 1470 5322 1504
rect 5356 1470 5399 1504
rect 5279 1430 5399 1470
rect 5279 1396 5322 1430
rect 5356 1396 5399 1430
rect 5279 1380 5399 1396
rect 5841 1504 5961 1552
rect 5841 1470 5884 1504
rect 5918 1470 5961 1504
rect 5841 1430 5961 1470
rect 5841 1396 5884 1430
rect 5918 1396 5961 1430
rect 5841 1380 5961 1396
rect 6271 1504 6391 1552
rect 6271 1470 6314 1504
rect 6348 1470 6391 1504
rect 6271 1430 6391 1470
rect 6271 1396 6314 1430
rect 6348 1396 6391 1430
rect 6271 1380 6391 1396
rect 6833 1504 6953 1552
rect 6833 1470 6876 1504
rect 6910 1470 6953 1504
rect 6833 1430 6953 1470
rect 6833 1396 6876 1430
rect 6910 1396 6953 1430
rect 6833 1380 6953 1396
rect 7263 1504 7383 1552
rect 7263 1470 7306 1504
rect 7340 1470 7383 1504
rect 7263 1430 7383 1470
rect 7263 1396 7306 1430
rect 7340 1396 7383 1430
rect 7263 1380 7383 1396
rect 7825 1504 7945 1552
rect 7825 1470 7868 1504
rect 7902 1470 7945 1504
rect 7825 1430 7945 1470
rect 7825 1396 7868 1430
rect 7902 1396 7945 1430
rect 7825 1380 7945 1396
rect 8255 1504 8375 1552
rect 8255 1470 8298 1504
rect 8332 1470 8375 1504
rect 8255 1430 8375 1470
rect 8255 1396 8298 1430
rect 8332 1396 8375 1430
rect 8255 1380 8375 1396
rect 8817 1504 8937 1552
rect 8817 1470 8860 1504
rect 8894 1470 8937 1504
rect 8817 1430 8937 1470
rect 8817 1396 8860 1430
rect 8894 1396 8937 1430
rect 8817 1380 8937 1396
rect 9247 1504 9367 1552
rect 9247 1470 9290 1504
rect 9324 1470 9367 1504
rect 9247 1430 9367 1470
rect 9247 1396 9290 1430
rect 9324 1396 9367 1430
rect 9247 1380 9367 1396
rect 9809 1504 9929 1552
rect 9809 1470 9852 1504
rect 9886 1470 9929 1504
rect 9809 1430 9929 1470
rect 9809 1396 9852 1430
rect 9886 1396 9929 1430
rect 9809 1380 9929 1396
rect 10239 1504 10359 1552
rect 10239 1470 10282 1504
rect 10316 1470 10359 1504
rect 10239 1430 10359 1470
rect 10239 1396 10282 1430
rect 10316 1396 10359 1430
rect 10239 1380 10359 1396
rect 10801 1504 10921 1552
rect 10801 1470 10844 1504
rect 10878 1470 10921 1504
rect 10801 1430 10921 1470
rect 10801 1396 10844 1430
rect 10878 1396 10921 1430
rect 10801 1380 10921 1396
rect 11231 1504 11351 1552
rect 11231 1470 11274 1504
rect 11308 1470 11351 1504
rect 11231 1430 11351 1470
rect 11231 1396 11274 1430
rect 11308 1396 11351 1430
rect 11231 1380 11351 1396
rect 11793 1504 11913 1552
rect 11793 1470 11836 1504
rect 11870 1470 11913 1504
rect 11793 1430 11913 1470
rect 11793 1396 11836 1430
rect 11870 1396 11913 1430
rect 11793 1380 11913 1396
rect 12223 1504 12343 1552
rect 12223 1470 12266 1504
rect 12300 1470 12343 1504
rect 12223 1430 12343 1470
rect 12223 1396 12266 1430
rect 12300 1396 12343 1430
rect 12223 1380 12343 1396
rect 12785 1504 12905 1552
rect 12785 1470 12828 1504
rect 12862 1470 12905 1504
rect 12785 1430 12905 1470
rect 12785 1396 12828 1430
rect 12862 1396 12905 1430
rect 12785 1380 12905 1396
rect 13215 1504 13335 1552
rect 13215 1470 13258 1504
rect 13292 1470 13335 1504
rect 13215 1430 13335 1470
rect 13215 1396 13258 1430
rect 13292 1396 13335 1430
rect 13215 1380 13335 1396
rect 13777 1504 13897 1552
rect 13777 1470 13820 1504
rect 13854 1470 13897 1504
rect 13777 1430 13897 1470
rect 13777 1396 13820 1430
rect 13854 1396 13897 1430
rect 13777 1380 13897 1396
rect 14135 1504 14255 1552
rect 14135 1470 14178 1504
rect 14212 1470 14255 1504
rect 14135 1430 14255 1470
rect 14135 1396 14178 1430
rect 14212 1396 14255 1430
rect 14135 1380 14255 1396
<< polycont >>
rect 924 4274 958 4308
rect 924 4200 958 4234
rect 1354 4274 1388 4308
rect 1354 4200 1388 4234
rect 1916 4274 1950 4308
rect 1916 4200 1950 4234
rect 2346 4274 2380 4308
rect 2346 4200 2380 4234
rect 2908 4274 2942 4308
rect 2908 4200 2942 4234
rect 3338 4274 3372 4308
rect 3338 4200 3372 4234
rect 3900 4274 3934 4308
rect 3900 4200 3934 4234
rect 4330 4274 4364 4308
rect 4330 4200 4364 4234
rect 4892 4274 4926 4308
rect 4892 4200 4926 4234
rect 5322 4274 5356 4308
rect 5322 4200 5356 4234
rect 5884 4274 5918 4308
rect 5884 4200 5918 4234
rect 6314 4274 6348 4308
rect 6314 4200 6348 4234
rect 6876 4274 6910 4308
rect 6876 4200 6910 4234
rect 7306 4274 7340 4308
rect 7306 4200 7340 4234
rect 7868 4274 7902 4308
rect 7868 4200 7902 4234
rect 8298 4274 8332 4308
rect 8298 4200 8332 4234
rect 8860 4274 8894 4308
rect 8860 4200 8894 4234
rect 9290 4274 9324 4308
rect 9290 4200 9324 4234
rect 9852 4274 9886 4308
rect 9852 4200 9886 4234
rect 10282 4274 10316 4308
rect 10282 4200 10316 4234
rect 10844 4274 10878 4308
rect 10844 4200 10878 4234
rect 11274 4274 11308 4308
rect 11274 4200 11308 4234
rect 11836 4274 11870 4308
rect 11836 4200 11870 4234
rect 12266 4274 12300 4308
rect 12266 4200 12300 4234
rect 12828 4274 12862 4308
rect 12828 4200 12862 4234
rect 13258 4274 13292 4308
rect 13258 4200 13292 4234
rect 13820 4274 13854 4308
rect 13820 4200 13854 4234
rect 14178 4274 14212 4308
rect 14178 4200 14212 4234
rect 924 3070 958 3104
rect 924 2992 958 3026
rect 924 2914 958 2948
rect 924 2836 958 2870
rect 924 2758 958 2792
rect 924 2679 958 2713
rect 924 2600 958 2634
rect 1354 3070 1388 3104
rect 1354 2992 1388 3026
rect 1354 2914 1388 2948
rect 1354 2836 1388 2870
rect 1354 2758 1388 2792
rect 1354 2679 1388 2713
rect 1354 2600 1388 2634
rect 1916 3070 1950 3104
rect 1916 2992 1950 3026
rect 1916 2914 1950 2948
rect 1916 2836 1950 2870
rect 1916 2758 1950 2792
rect 1916 2679 1950 2713
rect 1916 2600 1950 2634
rect 2346 3070 2380 3104
rect 2346 2992 2380 3026
rect 2346 2914 2380 2948
rect 2346 2836 2380 2870
rect 2346 2758 2380 2792
rect 2346 2679 2380 2713
rect 2346 2600 2380 2634
rect 2908 3070 2942 3104
rect 2908 2992 2942 3026
rect 2908 2914 2942 2948
rect 2908 2836 2942 2870
rect 2908 2758 2942 2792
rect 2908 2679 2942 2713
rect 2908 2600 2942 2634
rect 3338 3070 3372 3104
rect 3338 2992 3372 3026
rect 3338 2914 3372 2948
rect 3338 2836 3372 2870
rect 3338 2758 3372 2792
rect 3338 2679 3372 2713
rect 3338 2600 3372 2634
rect 3900 3070 3934 3104
rect 3900 2992 3934 3026
rect 3900 2914 3934 2948
rect 3900 2836 3934 2870
rect 3900 2758 3934 2792
rect 3900 2679 3934 2713
rect 3900 2600 3934 2634
rect 4330 3070 4364 3104
rect 4330 2992 4364 3026
rect 4330 2914 4364 2948
rect 4330 2836 4364 2870
rect 4330 2758 4364 2792
rect 4330 2679 4364 2713
rect 4330 2600 4364 2634
rect 4892 3070 4926 3104
rect 4892 2992 4926 3026
rect 4892 2914 4926 2948
rect 4892 2836 4926 2870
rect 4892 2758 4926 2792
rect 4892 2679 4926 2713
rect 4892 2600 4926 2634
rect 5322 3070 5356 3104
rect 5322 2992 5356 3026
rect 5322 2914 5356 2948
rect 5322 2836 5356 2870
rect 5322 2758 5356 2792
rect 5322 2679 5356 2713
rect 5322 2600 5356 2634
rect 5884 3070 5918 3104
rect 5884 2992 5918 3026
rect 5884 2914 5918 2948
rect 5884 2836 5918 2870
rect 5884 2758 5918 2792
rect 5884 2679 5918 2713
rect 5884 2600 5918 2634
rect 6314 3070 6348 3104
rect 6314 2992 6348 3026
rect 6314 2914 6348 2948
rect 6314 2836 6348 2870
rect 6314 2758 6348 2792
rect 6314 2679 6348 2713
rect 6314 2600 6348 2634
rect 6876 3070 6910 3104
rect 6876 2992 6910 3026
rect 6876 2914 6910 2948
rect 6876 2836 6910 2870
rect 6876 2758 6910 2792
rect 6876 2679 6910 2713
rect 6876 2600 6910 2634
rect 7306 3070 7340 3104
rect 7306 2992 7340 3026
rect 7306 2914 7340 2948
rect 7306 2836 7340 2870
rect 7306 2758 7340 2792
rect 7306 2679 7340 2713
rect 7306 2600 7340 2634
rect 7868 3070 7902 3104
rect 7868 2992 7902 3026
rect 7868 2914 7902 2948
rect 7868 2836 7902 2870
rect 7868 2758 7902 2792
rect 7868 2679 7902 2713
rect 7868 2600 7902 2634
rect 8298 3070 8332 3104
rect 8298 2992 8332 3026
rect 8298 2914 8332 2948
rect 8298 2836 8332 2870
rect 8298 2758 8332 2792
rect 8298 2679 8332 2713
rect 8298 2600 8332 2634
rect 8860 3070 8894 3104
rect 8860 2992 8894 3026
rect 8860 2914 8894 2948
rect 8860 2836 8894 2870
rect 8860 2758 8894 2792
rect 8860 2679 8894 2713
rect 8860 2600 8894 2634
rect 9290 3070 9324 3104
rect 9290 2992 9324 3026
rect 9290 2914 9324 2948
rect 9290 2836 9324 2870
rect 9290 2758 9324 2792
rect 9290 2679 9324 2713
rect 9290 2600 9324 2634
rect 9852 3070 9886 3104
rect 9852 2992 9886 3026
rect 9852 2914 9886 2948
rect 9852 2836 9886 2870
rect 9852 2758 9886 2792
rect 9852 2679 9886 2713
rect 9852 2600 9886 2634
rect 10282 3070 10316 3104
rect 10282 2992 10316 3026
rect 10282 2914 10316 2948
rect 10282 2836 10316 2870
rect 10282 2758 10316 2792
rect 10282 2679 10316 2713
rect 10282 2600 10316 2634
rect 10844 3070 10878 3104
rect 10844 2992 10878 3026
rect 10844 2914 10878 2948
rect 10844 2836 10878 2870
rect 10844 2758 10878 2792
rect 10844 2679 10878 2713
rect 10844 2600 10878 2634
rect 11274 3070 11308 3104
rect 11274 2992 11308 3026
rect 11274 2914 11308 2948
rect 11274 2836 11308 2870
rect 11274 2758 11308 2792
rect 11274 2679 11308 2713
rect 11274 2600 11308 2634
rect 11836 3070 11870 3104
rect 11836 2992 11870 3026
rect 11836 2914 11870 2948
rect 11836 2836 11870 2870
rect 11836 2758 11870 2792
rect 11836 2679 11870 2713
rect 11836 2600 11870 2634
rect 12266 3070 12300 3104
rect 12266 2992 12300 3026
rect 12266 2914 12300 2948
rect 12266 2836 12300 2870
rect 12266 2758 12300 2792
rect 12266 2679 12300 2713
rect 12266 2600 12300 2634
rect 12828 3070 12862 3104
rect 12828 2992 12862 3026
rect 12828 2914 12862 2948
rect 12828 2836 12862 2870
rect 12828 2758 12862 2792
rect 12828 2679 12862 2713
rect 12828 2600 12862 2634
rect 13258 3070 13292 3104
rect 13258 2992 13292 3026
rect 13258 2914 13292 2948
rect 13258 2836 13292 2870
rect 13258 2758 13292 2792
rect 13258 2679 13292 2713
rect 13258 2600 13292 2634
rect 13820 3070 13854 3104
rect 13820 2992 13854 3026
rect 13820 2914 13854 2948
rect 13820 2836 13854 2870
rect 13820 2758 13854 2792
rect 13820 2679 13854 2713
rect 13820 2600 13854 2634
rect 14178 3070 14212 3104
rect 14178 2992 14212 3026
rect 14178 2914 14212 2948
rect 14178 2836 14212 2870
rect 14178 2758 14212 2792
rect 14178 2679 14212 2713
rect 14178 2600 14212 2634
rect 924 1470 958 1504
rect 924 1396 958 1430
rect 1354 1470 1388 1504
rect 1354 1396 1388 1430
rect 1916 1470 1950 1504
rect 1916 1396 1950 1430
rect 2346 1470 2380 1504
rect 2346 1396 2380 1430
rect 2908 1470 2942 1504
rect 2908 1396 2942 1430
rect 3338 1470 3372 1504
rect 3338 1396 3372 1430
rect 3900 1470 3934 1504
rect 3900 1396 3934 1430
rect 4330 1470 4364 1504
rect 4330 1396 4364 1430
rect 4892 1470 4926 1504
rect 4892 1396 4926 1430
rect 5322 1470 5356 1504
rect 5322 1396 5356 1430
rect 5884 1470 5918 1504
rect 5884 1396 5918 1430
rect 6314 1470 6348 1504
rect 6314 1396 6348 1430
rect 6876 1470 6910 1504
rect 6876 1396 6910 1430
rect 7306 1470 7340 1504
rect 7306 1396 7340 1430
rect 7868 1470 7902 1504
rect 7868 1396 7902 1430
rect 8298 1470 8332 1504
rect 8298 1396 8332 1430
rect 8860 1470 8894 1504
rect 8860 1396 8894 1430
rect 9290 1470 9324 1504
rect 9290 1396 9324 1430
rect 9852 1470 9886 1504
rect 9852 1396 9886 1430
rect 10282 1470 10316 1504
rect 10282 1396 10316 1430
rect 10844 1470 10878 1504
rect 10844 1396 10878 1430
rect 11274 1470 11308 1504
rect 11274 1396 11308 1430
rect 11836 1470 11870 1504
rect 11836 1396 11870 1430
rect 12266 1470 12300 1504
rect 12266 1396 12300 1430
rect 12828 1470 12862 1504
rect 12828 1396 12862 1430
rect 13258 1470 13292 1504
rect 13258 1396 13292 1430
rect 13820 1470 13854 1504
rect 13820 1396 13854 1430
rect 14178 1470 14212 1504
rect 14178 1396 14212 1430
<< locali >>
rect 36 5111 15100 5118
rect 36 5077 361 5111
rect 395 5077 434 5111
rect 468 5077 507 5111
rect 541 5077 580 5111
rect 614 5077 653 5111
rect 687 5077 726 5111
rect 760 5077 799 5111
rect 833 5077 872 5111
rect 906 5077 945 5111
rect 979 5077 1018 5111
rect 1052 5077 1091 5111
rect 1125 5077 1164 5111
rect 1198 5077 1237 5111
rect 1271 5077 1310 5111
rect 1344 5077 1383 5111
rect 1417 5077 1456 5111
rect 1490 5077 1529 5111
rect 1563 5077 1602 5111
rect 1636 5077 1675 5111
rect 1709 5077 1748 5111
rect 1782 5077 1821 5111
rect 1855 5077 1894 5111
rect 1928 5077 1967 5111
rect 2001 5077 2040 5111
rect 2074 5077 2113 5111
rect 2147 5077 2186 5111
rect 2220 5077 2259 5111
rect 2293 5077 2332 5111
rect 2366 5077 2405 5111
rect 2439 5077 2478 5111
rect 2512 5077 2551 5111
rect 2585 5077 2624 5111
rect 2658 5077 2697 5111
rect 2731 5077 2770 5111
rect 2804 5077 2843 5111
rect 2877 5077 2916 5111
rect 2950 5077 2989 5111
rect 3023 5077 3062 5111
rect 3096 5077 3135 5111
rect 3169 5077 3208 5111
rect 3242 5077 3281 5111
rect 3315 5077 3354 5111
rect 3388 5077 3427 5111
rect 3461 5077 3500 5111
rect 3534 5077 3573 5111
rect 3607 5077 3646 5111
rect 3680 5077 3719 5111
rect 3753 5077 3792 5111
rect 3826 5077 3865 5111
rect 3899 5077 3938 5111
rect 3972 5077 4011 5111
rect 4045 5077 4084 5111
rect 4118 5077 4157 5111
rect 4191 5077 4229 5111
rect 4263 5077 4301 5111
rect 4335 5077 4373 5111
rect 4407 5077 4445 5111
rect 4479 5077 4517 5111
rect 4551 5077 4589 5111
rect 4623 5077 4661 5111
rect 4695 5077 4733 5111
rect 4767 5077 4805 5111
rect 4839 5077 4877 5111
rect 4911 5077 4949 5111
rect 4983 5077 5021 5111
rect 5055 5077 5093 5111
rect 5127 5077 5165 5111
rect 5199 5077 5237 5111
rect 5271 5077 5309 5111
rect 5343 5077 5381 5111
rect 5415 5077 5453 5111
rect 5487 5077 5525 5111
rect 5559 5077 5597 5111
rect 5631 5077 5669 5111
rect 5703 5077 5741 5111
rect 5775 5077 5813 5111
rect 5847 5077 5885 5111
rect 5919 5077 5957 5111
rect 5991 5077 6029 5111
rect 6063 5077 6101 5111
rect 6135 5077 6173 5111
rect 6207 5077 6245 5111
rect 6279 5077 6317 5111
rect 6351 5077 6389 5111
rect 6423 5077 6461 5111
rect 6495 5077 6533 5111
rect 6567 5077 6605 5111
rect 6639 5077 6677 5111
rect 6711 5077 6749 5111
rect 6783 5077 6821 5111
rect 6855 5077 6893 5111
rect 6927 5077 6965 5111
rect 6999 5077 7037 5111
rect 7071 5077 7109 5111
rect 7143 5077 7181 5111
rect 7215 5077 7253 5111
rect 7287 5077 7325 5111
rect 7359 5077 7397 5111
rect 7431 5077 7469 5111
rect 7503 5077 7541 5111
rect 7575 5077 7613 5111
rect 7647 5077 7685 5111
rect 7719 5077 7757 5111
rect 7791 5077 7829 5111
rect 7863 5077 7901 5111
rect 7935 5077 7973 5111
rect 8007 5077 8045 5111
rect 8079 5077 8117 5111
rect 8151 5077 8189 5111
rect 8223 5077 8261 5111
rect 8295 5077 8333 5111
rect 8367 5077 8405 5111
rect 8439 5077 8477 5111
rect 8511 5077 8549 5111
rect 8583 5077 8621 5111
rect 8655 5077 8693 5111
rect 8727 5077 8765 5111
rect 8799 5077 8837 5111
rect 8871 5077 8909 5111
rect 8943 5077 8981 5111
rect 9015 5077 9053 5111
rect 9087 5077 9125 5111
rect 9159 5077 9197 5111
rect 9231 5077 9269 5111
rect 9303 5077 9341 5111
rect 9375 5077 9413 5111
rect 9447 5077 9485 5111
rect 9519 5077 9557 5111
rect 9591 5077 9629 5111
rect 9663 5077 9701 5111
rect 9735 5077 9773 5111
rect 9807 5077 9845 5111
rect 9879 5077 9917 5111
rect 9951 5077 9989 5111
rect 10023 5077 10061 5111
rect 10095 5077 10133 5111
rect 10167 5077 10205 5111
rect 10239 5077 10277 5111
rect 10311 5077 10349 5111
rect 10383 5077 10421 5111
rect 10455 5077 10493 5111
rect 10527 5077 10565 5111
rect 10599 5077 10637 5111
rect 10671 5077 10709 5111
rect 10743 5077 10781 5111
rect 10815 5077 10853 5111
rect 10887 5077 10925 5111
rect 10959 5077 10997 5111
rect 11031 5077 11069 5111
rect 11103 5077 11141 5111
rect 11175 5077 11213 5111
rect 11247 5077 11285 5111
rect 11319 5077 11357 5111
rect 11391 5077 11429 5111
rect 11463 5077 11501 5111
rect 11535 5077 11573 5111
rect 11607 5077 11645 5111
rect 11679 5077 11717 5111
rect 11751 5077 11789 5111
rect 11823 5077 11861 5111
rect 11895 5077 11933 5111
rect 11967 5077 12005 5111
rect 12039 5077 12077 5111
rect 12111 5077 12149 5111
rect 12183 5077 12221 5111
rect 12255 5077 12293 5111
rect 12327 5077 12365 5111
rect 12399 5077 12437 5111
rect 12471 5077 12509 5111
rect 12543 5077 12581 5111
rect 12615 5077 12653 5111
rect 12687 5077 12725 5111
rect 12759 5077 12797 5111
rect 12831 5077 12869 5111
rect 12903 5077 12941 5111
rect 12975 5077 13013 5111
rect 13047 5077 13085 5111
rect 13119 5077 13157 5111
rect 13191 5077 13229 5111
rect 13263 5077 13301 5111
rect 13335 5077 13373 5111
rect 13407 5077 13445 5111
rect 13479 5077 13517 5111
rect 13551 5077 13589 5111
rect 13623 5077 13661 5111
rect 13695 5077 13733 5111
rect 13767 5077 13805 5111
rect 13839 5077 13877 5111
rect 13911 5077 13949 5111
rect 13983 5077 14021 5111
rect 14055 5077 14093 5111
rect 14127 5077 14165 5111
rect 14199 5077 14237 5111
rect 14271 5077 14309 5111
rect 14343 5077 14381 5111
rect 14415 5077 14453 5111
rect 14487 5077 14525 5111
rect 14559 5077 14597 5111
rect 14631 5077 14669 5111
rect 14703 5077 14741 5111
rect 14775 5077 15100 5111
rect 36 5068 15100 5077
rect 36 5049 142 5068
rect 36 331 51 5049
rect 85 5045 142 5049
rect 176 5045 214 5068
rect 248 5034 286 5068
rect 320 5034 358 5068
rect 392 5035 430 5068
rect 464 5035 502 5068
rect 536 5035 574 5068
rect 608 5035 646 5068
rect 680 5035 718 5068
rect 752 5035 790 5068
rect 824 5035 862 5068
rect 896 5035 934 5068
rect 968 5035 1006 5068
rect 1040 5035 1078 5068
rect 1112 5035 1150 5068
rect 1184 5035 1222 5068
rect 1256 5035 1294 5068
rect 1328 5035 1366 5068
rect 1400 5035 1438 5068
rect 1472 5035 1510 5068
rect 1544 5035 1582 5068
rect 1616 5035 1654 5068
rect 1688 5035 1726 5068
rect 1760 5035 1798 5068
rect 1832 5035 1870 5068
rect 1904 5035 1942 5068
rect 1976 5035 2014 5068
rect 2048 5035 2086 5068
rect 2120 5035 2158 5068
rect 2192 5035 2230 5068
rect 2264 5035 2302 5068
rect 2336 5035 2374 5068
rect 2408 5035 2446 5068
rect 2480 5035 2518 5068
rect 2552 5035 2590 5068
rect 395 5034 430 5035
rect 468 5034 502 5035
rect 541 5034 574 5035
rect 614 5034 646 5035
rect 687 5034 718 5035
rect 760 5034 790 5035
rect 833 5034 862 5035
rect 906 5034 934 5035
rect 979 5034 1006 5035
rect 1052 5034 1078 5035
rect 1125 5034 1150 5035
rect 1198 5034 1222 5035
rect 1271 5034 1294 5035
rect 1344 5034 1366 5035
rect 1417 5034 1438 5035
rect 1490 5034 1510 5035
rect 1563 5034 1582 5035
rect 1636 5034 1654 5035
rect 1709 5034 1726 5035
rect 1782 5034 1798 5035
rect 1855 5034 1870 5035
rect 1928 5034 1942 5035
rect 2001 5034 2014 5035
rect 2074 5034 2086 5035
rect 2147 5034 2158 5035
rect 2220 5034 2230 5035
rect 2293 5034 2302 5035
rect 2366 5034 2374 5035
rect 2439 5034 2446 5035
rect 2512 5034 2518 5035
rect 2585 5034 2590 5035
rect 2624 5035 2662 5068
rect 229 5029 361 5034
rect 229 5000 269 5029
rect 303 5001 361 5029
rect 395 5001 434 5034
rect 468 5001 507 5034
rect 541 5001 580 5034
rect 614 5001 653 5034
rect 687 5001 726 5034
rect 760 5001 799 5034
rect 833 5001 872 5034
rect 906 5001 945 5034
rect 979 5001 1018 5034
rect 1052 5001 1091 5034
rect 1125 5001 1164 5034
rect 1198 5001 1237 5034
rect 1271 5001 1310 5034
rect 1344 5001 1383 5034
rect 1417 5001 1456 5034
rect 1490 5001 1529 5034
rect 1563 5001 1602 5034
rect 1636 5001 1675 5034
rect 1709 5001 1748 5034
rect 1782 5001 1821 5034
rect 1855 5001 1894 5034
rect 1928 5001 1967 5034
rect 2001 5001 2040 5034
rect 2074 5001 2113 5034
rect 2147 5001 2186 5034
rect 2220 5001 2259 5034
rect 2293 5001 2332 5034
rect 2366 5001 2405 5034
rect 2439 5001 2478 5034
rect 2512 5001 2551 5034
rect 2585 5001 2624 5034
rect 2658 5034 2662 5035
rect 2696 5035 2734 5068
rect 2696 5034 2697 5035
rect 2658 5001 2697 5034
rect 2731 5034 2734 5035
rect 2768 5035 2806 5068
rect 2768 5034 2770 5035
rect 2731 5001 2770 5034
rect 2804 5034 2806 5035
rect 2840 5035 2878 5068
rect 2840 5034 2843 5035
rect 2804 5001 2843 5034
rect 2877 5034 2878 5035
rect 2912 5035 2950 5068
rect 2912 5034 2916 5035
rect 2877 5001 2916 5034
rect 2984 5035 3022 5068
rect 3056 5035 3094 5068
rect 3128 5035 3166 5068
rect 3200 5035 3238 5068
rect 3272 5035 3310 5068
rect 3344 5035 3382 5068
rect 3416 5035 3454 5068
rect 3488 5035 3526 5068
rect 3560 5035 3598 5068
rect 3632 5035 3670 5068
rect 3704 5035 3742 5068
rect 3776 5035 3814 5068
rect 3848 5035 3886 5068
rect 3920 5035 3958 5068
rect 3992 5035 4030 5068
rect 4064 5035 4102 5068
rect 4136 5035 4174 5068
rect 4208 5035 4246 5068
rect 4280 5035 4318 5068
rect 4352 5035 4390 5068
rect 4424 5035 4462 5068
rect 4496 5035 4534 5068
rect 4568 5035 4606 5068
rect 4640 5035 4678 5068
rect 4712 5035 4750 5068
rect 4784 5035 4822 5068
rect 4856 5035 4894 5068
rect 4928 5035 4966 5068
rect 5000 5035 5038 5068
rect 5072 5035 5110 5068
rect 5144 5035 5182 5068
rect 5216 5035 5254 5068
rect 5288 5035 5326 5068
rect 5360 5035 5398 5068
rect 5432 5035 5470 5068
rect 5504 5035 5542 5068
rect 5576 5035 5614 5068
rect 5648 5035 5686 5068
rect 5720 5035 5758 5068
rect 5792 5035 5830 5068
rect 5864 5035 5902 5068
rect 5936 5035 5974 5068
rect 6008 5035 6046 5068
rect 6080 5035 6118 5068
rect 6152 5035 6190 5068
rect 6224 5035 6262 5068
rect 6296 5035 6334 5068
rect 6368 5035 6406 5068
rect 6440 5035 6478 5068
rect 6512 5035 6550 5068
rect 6584 5035 6622 5068
rect 6656 5035 6694 5068
rect 6728 5035 6766 5068
rect 6800 5035 6838 5068
rect 6872 5035 6910 5068
rect 6944 5035 6982 5068
rect 7016 5035 7054 5068
rect 7088 5035 7126 5068
rect 7160 5035 7198 5068
rect 7232 5035 7270 5068
rect 7304 5035 7342 5068
rect 7376 5035 7414 5068
rect 7448 5035 7486 5068
rect 7520 5035 7558 5068
rect 7592 5035 7630 5068
rect 7664 5035 7702 5068
rect 7736 5035 7774 5068
rect 7808 5035 7846 5068
rect 7880 5035 7918 5068
rect 7952 5035 7990 5068
rect 8024 5035 8062 5068
rect 8096 5035 8134 5068
rect 8168 5035 8206 5068
rect 8240 5035 8278 5068
rect 8312 5035 8350 5068
rect 8384 5035 8422 5068
rect 8456 5035 8494 5068
rect 8528 5035 8566 5068
rect 8600 5035 8638 5068
rect 8672 5035 8710 5068
rect 8744 5035 8782 5068
rect 8816 5035 8854 5068
rect 8888 5035 8926 5068
rect 8960 5035 8998 5068
rect 9032 5035 9070 5068
rect 9104 5035 9142 5068
rect 9176 5035 9214 5068
rect 9248 5035 9286 5068
rect 9320 5035 9358 5068
rect 9392 5035 9430 5068
rect 9464 5035 9502 5068
rect 9536 5035 9574 5068
rect 9608 5035 9646 5068
rect 9680 5035 9718 5068
rect 9752 5035 9790 5068
rect 9824 5035 9862 5068
rect 9896 5035 9934 5068
rect 9968 5035 10006 5068
rect 10040 5035 10078 5068
rect 10112 5035 10151 5068
rect 10185 5035 10224 5068
rect 10258 5035 10297 5068
rect 10331 5035 10370 5068
rect 10404 5035 10443 5068
rect 10477 5035 10516 5068
rect 10550 5035 10589 5068
rect 10623 5035 10662 5068
rect 10696 5035 10735 5068
rect 10769 5035 10808 5068
rect 10842 5035 10881 5068
rect 10915 5035 10954 5068
rect 10988 5035 11027 5068
rect 11061 5035 11100 5068
rect 11134 5035 11173 5068
rect 11207 5035 11246 5068
rect 11280 5035 11319 5068
rect 2984 5034 2989 5035
rect 3056 5034 3062 5035
rect 3128 5034 3135 5035
rect 3200 5034 3208 5035
rect 3272 5034 3281 5035
rect 3344 5034 3354 5035
rect 3416 5034 3427 5035
rect 3488 5034 3500 5035
rect 3560 5034 3573 5035
rect 3632 5034 3646 5035
rect 3704 5034 3719 5035
rect 3776 5034 3792 5035
rect 3848 5034 3865 5035
rect 3920 5034 3938 5035
rect 3992 5034 4011 5035
rect 4064 5034 4084 5035
rect 4136 5034 4157 5035
rect 4208 5034 4229 5035
rect 4280 5034 4301 5035
rect 4352 5034 4373 5035
rect 4424 5034 4445 5035
rect 4496 5034 4517 5035
rect 4568 5034 4589 5035
rect 4640 5034 4661 5035
rect 4712 5034 4733 5035
rect 4784 5034 4805 5035
rect 4856 5034 4877 5035
rect 4928 5034 4949 5035
rect 5000 5034 5021 5035
rect 5072 5034 5093 5035
rect 5144 5034 5165 5035
rect 5216 5034 5237 5035
rect 5288 5034 5309 5035
rect 5360 5034 5381 5035
rect 5432 5034 5453 5035
rect 5504 5034 5525 5035
rect 5576 5034 5597 5035
rect 5648 5034 5669 5035
rect 5720 5034 5741 5035
rect 5792 5034 5813 5035
rect 5864 5034 5885 5035
rect 5936 5034 5957 5035
rect 6008 5034 6029 5035
rect 6080 5034 6101 5035
rect 6152 5034 6173 5035
rect 6224 5034 6245 5035
rect 6296 5034 6317 5035
rect 6368 5034 6389 5035
rect 6440 5034 6461 5035
rect 6512 5034 6533 5035
rect 6584 5034 6605 5035
rect 6656 5034 6677 5035
rect 6728 5034 6749 5035
rect 6800 5034 6821 5035
rect 6872 5034 6893 5035
rect 6944 5034 6965 5035
rect 7016 5034 7037 5035
rect 7088 5034 7109 5035
rect 7160 5034 7181 5035
rect 7232 5034 7253 5035
rect 7304 5034 7325 5035
rect 7376 5034 7397 5035
rect 7448 5034 7469 5035
rect 7520 5034 7541 5035
rect 7592 5034 7613 5035
rect 7664 5034 7685 5035
rect 7736 5034 7757 5035
rect 7808 5034 7829 5035
rect 7880 5034 7901 5035
rect 7952 5034 7973 5035
rect 8024 5034 8045 5035
rect 8096 5034 8117 5035
rect 8168 5034 8189 5035
rect 8240 5034 8261 5035
rect 8312 5034 8333 5035
rect 8384 5034 8405 5035
rect 8456 5034 8477 5035
rect 8528 5034 8549 5035
rect 8600 5034 8621 5035
rect 8672 5034 8693 5035
rect 8744 5034 8765 5035
rect 8816 5034 8837 5035
rect 8888 5034 8909 5035
rect 8960 5034 8981 5035
rect 9032 5034 9053 5035
rect 9104 5034 9125 5035
rect 9176 5034 9197 5035
rect 9248 5034 9269 5035
rect 9320 5034 9341 5035
rect 9392 5034 9413 5035
rect 9464 5034 9485 5035
rect 9536 5034 9557 5035
rect 9608 5034 9629 5035
rect 9680 5034 9701 5035
rect 9752 5034 9773 5035
rect 9824 5034 9845 5035
rect 9896 5034 9917 5035
rect 9968 5034 9989 5035
rect 10040 5034 10061 5035
rect 10112 5034 10133 5035
rect 10185 5034 10205 5035
rect 10258 5034 10277 5035
rect 10331 5034 10349 5035
rect 10404 5034 10421 5035
rect 10477 5034 10493 5035
rect 10550 5034 10565 5035
rect 10623 5034 10637 5035
rect 10696 5034 10709 5035
rect 10769 5034 10781 5035
rect 10842 5034 10853 5035
rect 10915 5034 10925 5035
rect 10988 5034 10997 5035
rect 11061 5034 11069 5035
rect 11134 5034 11141 5035
rect 11207 5034 11213 5035
rect 11280 5034 11285 5035
rect 2950 5001 2989 5034
rect 3023 5001 3062 5034
rect 3096 5001 3135 5034
rect 3169 5001 3208 5034
rect 3242 5001 3281 5034
rect 3315 5001 3354 5034
rect 3388 5001 3427 5034
rect 3461 5001 3500 5034
rect 3534 5001 3573 5034
rect 3607 5001 3646 5034
rect 3680 5001 3719 5034
rect 3753 5001 3792 5034
rect 3826 5001 3865 5034
rect 3899 5001 3938 5034
rect 3972 5001 4011 5034
rect 4045 5001 4084 5034
rect 4118 5001 4157 5034
rect 4191 5001 4229 5034
rect 4263 5001 4301 5034
rect 4335 5001 4373 5034
rect 4407 5001 4445 5034
rect 4479 5001 4517 5034
rect 4551 5001 4589 5034
rect 4623 5001 4661 5034
rect 4695 5001 4733 5034
rect 4767 5001 4805 5034
rect 4839 5001 4877 5034
rect 4911 5001 4949 5034
rect 4983 5001 5021 5034
rect 5055 5001 5093 5034
rect 5127 5001 5165 5034
rect 5199 5001 5237 5034
rect 5271 5001 5309 5034
rect 5343 5001 5381 5034
rect 5415 5001 5453 5034
rect 5487 5001 5525 5034
rect 5559 5001 5597 5034
rect 5631 5001 5669 5034
rect 5703 5001 5741 5034
rect 5775 5001 5813 5034
rect 5847 5001 5885 5034
rect 5919 5001 5957 5034
rect 5991 5001 6029 5034
rect 6063 5001 6101 5034
rect 6135 5001 6173 5034
rect 6207 5001 6245 5034
rect 6279 5001 6317 5034
rect 6351 5001 6389 5034
rect 6423 5001 6461 5034
rect 6495 5001 6533 5034
rect 6567 5001 6605 5034
rect 6639 5001 6677 5034
rect 6711 5001 6749 5034
rect 6783 5001 6821 5034
rect 6855 5001 6893 5034
rect 6927 5001 6965 5034
rect 6999 5001 7037 5034
rect 7071 5001 7109 5034
rect 7143 5001 7181 5034
rect 7215 5001 7253 5034
rect 7287 5001 7325 5034
rect 7359 5001 7397 5034
rect 7431 5001 7469 5034
rect 7503 5001 7541 5034
rect 7575 5001 7613 5034
rect 7647 5001 7685 5034
rect 7719 5001 7757 5034
rect 7791 5001 7829 5034
rect 7863 5001 7901 5034
rect 7935 5001 7973 5034
rect 8007 5001 8045 5034
rect 8079 5001 8117 5034
rect 8151 5001 8189 5034
rect 8223 5001 8261 5034
rect 8295 5001 8333 5034
rect 8367 5001 8405 5034
rect 8439 5001 8477 5034
rect 8511 5001 8549 5034
rect 8583 5001 8621 5034
rect 8655 5001 8693 5034
rect 8727 5001 8765 5034
rect 8799 5001 8837 5034
rect 8871 5001 8909 5034
rect 8943 5001 8981 5034
rect 9015 5001 9053 5034
rect 9087 5001 9125 5034
rect 9159 5001 9197 5034
rect 9231 5001 9269 5034
rect 9303 5001 9341 5034
rect 9375 5001 9413 5034
rect 9447 5001 9485 5034
rect 9519 5001 9557 5034
rect 9591 5001 9629 5034
rect 9663 5001 9701 5034
rect 9735 5001 9773 5034
rect 9807 5001 9845 5034
rect 9879 5001 9917 5034
rect 9951 5001 9989 5034
rect 10023 5001 10061 5034
rect 10095 5001 10133 5034
rect 10167 5001 10205 5034
rect 10239 5001 10277 5034
rect 10311 5001 10349 5034
rect 10383 5001 10421 5034
rect 10455 5001 10493 5034
rect 10527 5001 10565 5034
rect 10599 5001 10637 5034
rect 10671 5001 10709 5034
rect 10743 5001 10781 5034
rect 10815 5001 10853 5034
rect 10887 5001 10925 5034
rect 10959 5001 10997 5034
rect 11031 5001 11069 5034
rect 11103 5001 11141 5034
rect 11175 5001 11213 5034
rect 11247 5001 11285 5034
rect 11353 5035 11392 5068
rect 11353 5034 11357 5035
rect 11319 5001 11357 5034
rect 11391 5034 11392 5035
rect 11426 5035 11465 5068
rect 11426 5034 11429 5035
rect 11391 5001 11429 5034
rect 11463 5034 11465 5035
rect 11499 5035 11538 5068
rect 11499 5034 11501 5035
rect 11463 5001 11501 5034
rect 11535 5034 11538 5035
rect 11572 5035 11611 5068
rect 11572 5034 11573 5035
rect 11535 5001 11573 5034
rect 11607 5034 11611 5035
rect 11645 5035 11684 5068
rect 11718 5035 11757 5068
rect 11791 5035 11830 5068
rect 11864 5035 11903 5068
rect 11937 5035 11976 5068
rect 12010 5035 12049 5068
rect 12083 5035 12122 5068
rect 12156 5035 12195 5068
rect 12229 5035 12268 5068
rect 12302 5035 12341 5068
rect 12375 5035 12414 5068
rect 12448 5035 12487 5068
rect 12521 5035 12560 5068
rect 12594 5035 12633 5068
rect 12667 5035 12706 5068
rect 12740 5035 12779 5068
rect 12813 5035 12852 5068
rect 12886 5035 12925 5068
rect 12959 5035 12998 5068
rect 13032 5035 13071 5068
rect 13105 5035 13144 5068
rect 13178 5035 13217 5068
rect 13251 5035 13290 5068
rect 13324 5035 13363 5068
rect 13397 5035 13436 5068
rect 13470 5035 13509 5068
rect 13543 5035 13582 5068
rect 13616 5035 13655 5068
rect 13689 5035 13728 5068
rect 13762 5035 13801 5068
rect 13835 5035 13874 5068
rect 13908 5035 13947 5068
rect 13981 5035 14020 5068
rect 14054 5035 14093 5068
rect 14127 5035 14166 5068
rect 14200 5035 14239 5068
rect 14273 5035 14312 5068
rect 14346 5035 14385 5068
rect 14419 5035 14458 5068
rect 14492 5035 14531 5068
rect 14565 5035 14604 5068
rect 14638 5035 14677 5068
rect 14711 5035 14750 5068
rect 11607 5001 11645 5034
rect 11679 5034 11684 5035
rect 11751 5034 11757 5035
rect 11823 5034 11830 5035
rect 11895 5034 11903 5035
rect 11967 5034 11976 5035
rect 12039 5034 12049 5035
rect 12111 5034 12122 5035
rect 12183 5034 12195 5035
rect 12255 5034 12268 5035
rect 12327 5034 12341 5035
rect 12399 5034 12414 5035
rect 12471 5034 12487 5035
rect 12543 5034 12560 5035
rect 12615 5034 12633 5035
rect 12687 5034 12706 5035
rect 12759 5034 12779 5035
rect 12831 5034 12852 5035
rect 12903 5034 12925 5035
rect 12975 5034 12998 5035
rect 13047 5034 13071 5035
rect 13119 5034 13144 5035
rect 13191 5034 13217 5035
rect 13263 5034 13290 5035
rect 13335 5034 13363 5035
rect 13407 5034 13436 5035
rect 13479 5034 13509 5035
rect 13551 5034 13582 5035
rect 13623 5034 13655 5035
rect 13695 5034 13728 5035
rect 13767 5034 13801 5035
rect 13839 5034 13874 5035
rect 13911 5034 13947 5035
rect 13983 5034 14020 5035
rect 11679 5001 11717 5034
rect 11751 5001 11789 5034
rect 11823 5001 11861 5034
rect 11895 5001 11933 5034
rect 11967 5001 12005 5034
rect 12039 5001 12077 5034
rect 12111 5001 12149 5034
rect 12183 5001 12221 5034
rect 12255 5001 12293 5034
rect 12327 5001 12365 5034
rect 12399 5001 12437 5034
rect 12471 5001 12509 5034
rect 12543 5001 12581 5034
rect 12615 5001 12653 5034
rect 12687 5001 12725 5034
rect 12759 5001 12797 5034
rect 12831 5001 12869 5034
rect 12903 5001 12941 5034
rect 12975 5001 13013 5034
rect 13047 5001 13085 5034
rect 13119 5001 13157 5034
rect 13191 5001 13229 5034
rect 13263 5001 13301 5034
rect 13335 5001 13373 5034
rect 13407 5001 13445 5034
rect 13479 5001 13517 5034
rect 13551 5001 13589 5034
rect 13623 5001 13661 5034
rect 13695 5001 13733 5034
rect 13767 5001 13805 5034
rect 13839 5001 13877 5034
rect 13911 5001 13949 5034
rect 13983 5001 14021 5034
rect 14055 5001 14093 5035
rect 14127 5001 14165 5035
rect 14200 5034 14237 5035
rect 14273 5034 14309 5035
rect 14346 5034 14381 5035
rect 14419 5034 14453 5035
rect 14492 5034 14525 5035
rect 14565 5034 14597 5035
rect 14638 5034 14669 5035
rect 14711 5034 14741 5035
rect 14784 5034 14823 5068
rect 14857 5062 15100 5068
rect 14857 5034 14907 5062
rect 14199 5001 14237 5034
rect 14271 5001 14309 5034
rect 14343 5001 14381 5034
rect 14415 5001 14453 5034
rect 14487 5001 14525 5034
rect 14559 5001 14597 5034
rect 14631 5001 14669 5034
rect 14703 5001 14741 5034
rect 14775 5030 14907 5034
rect 14775 5001 14832 5030
rect 303 5000 14832 5001
rect 229 4966 263 5000
rect 303 4995 335 5000
rect 297 4966 335 4995
rect 369 4966 407 5000
rect 441 4966 479 5000
rect 513 4966 551 5000
rect 585 4966 623 5000
rect 657 4966 695 5000
rect 729 4966 767 5000
rect 801 4966 839 5000
rect 873 4966 911 5000
rect 945 4966 983 5000
rect 1017 4966 1055 5000
rect 1089 4966 1127 5000
rect 1161 4966 1199 5000
rect 1233 4966 1271 5000
rect 1305 4966 1343 5000
rect 1377 4966 1415 5000
rect 1449 4966 1487 5000
rect 1521 4966 1559 5000
rect 1593 4966 1631 5000
rect 1665 4966 1703 5000
rect 1737 4966 1775 5000
rect 1809 4966 1847 5000
rect 1881 4966 1919 5000
rect 1953 4966 1991 5000
rect 2025 4966 2063 5000
rect 2097 4966 2135 5000
rect 2169 4966 2207 5000
rect 2241 4966 2279 5000
rect 2313 4966 2351 5000
rect 2385 4966 2423 5000
rect 2457 4966 2495 5000
rect 2529 4966 2567 5000
rect 2601 4966 2639 5000
rect 2673 4966 2711 5000
rect 2745 4966 2783 5000
rect 2817 4966 2855 5000
rect 2889 4966 2927 5000
rect 2961 4966 2999 5000
rect 3033 4966 3071 5000
rect 3105 4966 3143 5000
rect 3177 4966 3215 5000
rect 3249 4966 3287 5000
rect 3321 4966 3359 5000
rect 3393 4966 3431 5000
rect 3465 4966 3503 5000
rect 3537 4966 3575 5000
rect 3609 4966 3647 5000
rect 3681 4966 3719 5000
rect 3753 4966 3791 5000
rect 3825 4966 3863 5000
rect 3897 4966 3935 5000
rect 3969 4966 4007 5000
rect 4041 4966 4079 5000
rect 4113 4966 4151 5000
rect 4185 4966 4223 5000
rect 4257 4966 4295 5000
rect 4329 4966 4367 5000
rect 4401 4966 4439 5000
rect 4473 4966 4511 5000
rect 4545 4966 4583 5000
rect 4617 4966 4655 5000
rect 4689 4966 4727 5000
rect 4761 4966 4799 5000
rect 4833 4966 4871 5000
rect 4905 4966 4943 5000
rect 4977 4966 5015 5000
rect 5049 4966 5087 5000
rect 5121 4966 5159 5000
rect 5193 4966 5231 5000
rect 5265 4966 5303 5000
rect 5337 4966 5375 5000
rect 5409 4966 5447 5000
rect 5481 4966 5519 5000
rect 5553 4966 5591 5000
rect 5625 4966 5663 5000
rect 5697 4966 5735 5000
rect 5769 4966 5807 5000
rect 5841 4966 5879 5000
rect 5913 4966 5951 5000
rect 5985 4966 6023 5000
rect 6057 4966 6095 5000
rect 6129 4966 6167 5000
rect 6201 4966 6239 5000
rect 6273 4966 6311 5000
rect 6345 4966 6383 5000
rect 6417 4966 6455 5000
rect 6489 4966 6527 5000
rect 6561 4966 6599 5000
rect 6633 4966 6671 5000
rect 6705 4966 6743 5000
rect 6777 4966 6815 5000
rect 6849 4966 6887 5000
rect 6921 4966 6959 5000
rect 6993 4966 7031 5000
rect 7065 4966 7103 5000
rect 7137 4966 7175 5000
rect 7209 4966 7247 5000
rect 7281 4966 7319 5000
rect 7353 4966 7391 5000
rect 7425 4966 7463 5000
rect 7497 4966 7535 5000
rect 7569 4966 7607 5000
rect 7641 4966 7679 5000
rect 7713 4966 7751 5000
rect 7785 4966 7823 5000
rect 7857 4966 7895 5000
rect 7929 4966 7967 5000
rect 8001 4966 8039 5000
rect 8073 4966 8111 5000
rect 8145 4966 8183 5000
rect 8217 4966 8255 5000
rect 8289 4966 8327 5000
rect 8361 4966 8399 5000
rect 8433 4966 8471 5000
rect 8505 4966 8543 5000
rect 8577 4966 8615 5000
rect 8649 4966 8687 5000
rect 8721 4966 8759 5000
rect 8793 4966 8831 5000
rect 8865 4966 8903 5000
rect 8937 4966 8975 5000
rect 9009 4966 9047 5000
rect 9081 4966 9119 5000
rect 9153 4966 9191 5000
rect 9225 4966 9263 5000
rect 9297 4966 9335 5000
rect 9369 4966 9407 5000
rect 9441 4966 9479 5000
rect 9513 4966 9551 5000
rect 9585 4966 9623 5000
rect 9657 4966 9695 5000
rect 9729 4966 9767 5000
rect 9801 4966 9839 5000
rect 9873 4966 9911 5000
rect 9945 4966 9983 5000
rect 10017 4966 10055 5000
rect 10089 4966 10127 5000
rect 10161 4966 10199 5000
rect 10233 4966 10271 5000
rect 10305 4966 10343 5000
rect 10377 4966 10415 5000
rect 10449 4966 10487 5000
rect 10521 4966 10559 5000
rect 10593 4966 10631 5000
rect 10665 4966 10703 5000
rect 10737 4966 10775 5000
rect 10809 4966 10847 5000
rect 10881 4966 10919 5000
rect 10953 4966 10991 5000
rect 11025 4966 11063 5000
rect 11097 4966 11135 5000
rect 11169 4966 11207 5000
rect 11241 4966 11279 5000
rect 11313 4966 11351 5000
rect 11385 4966 11423 5000
rect 11457 4966 11495 5000
rect 11529 4966 11567 5000
rect 11601 4966 11639 5000
rect 11673 4966 11711 5000
rect 11745 4966 11783 5000
rect 11817 4966 11855 5000
rect 11889 4966 11927 5000
rect 11961 4966 11999 5000
rect 12033 4966 12071 5000
rect 12105 4966 12143 5000
rect 12177 4966 12215 5000
rect 12249 4966 12287 5000
rect 12321 4966 12359 5000
rect 12393 4966 12431 5000
rect 12465 4966 12503 5000
rect 12537 4966 12575 5000
rect 12609 4966 12647 5000
rect 12681 4966 12719 5000
rect 12753 4966 12791 5000
rect 12825 4966 12863 5000
rect 12897 4966 12935 5000
rect 12969 4966 13007 5000
rect 13041 4966 13079 5000
rect 13113 4966 13151 5000
rect 13185 4966 13223 5000
rect 13257 4966 13295 5000
rect 13329 4966 13367 5000
rect 13401 4966 13439 5000
rect 13473 4966 13511 5000
rect 13545 4966 13583 5000
rect 13617 4966 13655 5000
rect 13689 4966 13728 5000
rect 13762 4966 13801 5000
rect 13835 4966 13874 5000
rect 13908 4966 13947 5000
rect 13981 4966 14020 5000
rect 14054 4966 14093 5000
rect 14127 4966 14166 5000
rect 14200 4966 14239 5000
rect 14273 4966 14312 5000
rect 14346 4966 14385 5000
rect 14419 4966 14458 5000
rect 14492 4966 14531 5000
rect 14565 4966 14604 5000
rect 14638 4966 14677 5000
rect 14711 4966 14750 5000
rect 14784 4966 14823 5000
rect 14866 4996 14907 5030
rect 14857 4966 14907 4996
rect 229 4959 14907 4966
rect 229 4956 361 4959
rect 229 4932 269 4956
rect 303 4932 361 4956
rect 395 4932 434 4959
rect 468 4932 507 4959
rect 541 4932 580 4959
rect 614 4932 653 4959
rect 229 4898 259 4932
rect 303 4922 331 4932
rect 395 4925 403 4932
rect 468 4925 475 4932
rect 541 4925 547 4932
rect 614 4925 619 4932
rect 293 4898 331 4922
rect 365 4898 403 4925
rect 437 4898 475 4925
rect 509 4898 547 4925
rect 581 4898 619 4925
rect 687 4932 726 4959
rect 687 4925 691 4932
rect 653 4898 691 4925
rect 725 4925 726 4932
rect 760 4932 799 4959
rect 760 4925 763 4932
rect 725 4898 763 4925
rect 797 4925 799 4932
rect 833 4932 872 4959
rect 833 4925 835 4932
rect 797 4898 835 4925
rect 869 4925 872 4932
rect 906 4932 945 4959
rect 906 4925 907 4932
rect 869 4898 907 4925
rect 941 4925 945 4932
rect 979 4932 1018 4959
rect 1052 4932 1091 4959
rect 1125 4932 1164 4959
rect 1198 4932 1237 4959
rect 1271 4932 1310 4959
rect 1344 4932 1383 4959
rect 1417 4932 1456 4959
rect 1490 4932 1529 4959
rect 1563 4932 1602 4959
rect 1636 4932 1675 4959
rect 1709 4932 1748 4959
rect 1782 4932 1821 4959
rect 1855 4932 1894 4959
rect 1928 4932 1967 4959
rect 2001 4932 2040 4959
rect 2074 4932 2113 4959
rect 2147 4932 2186 4959
rect 2220 4932 2259 4959
rect 2293 4932 2332 4959
rect 2366 4932 2405 4959
rect 2439 4932 2478 4959
rect 2512 4932 2551 4959
rect 2585 4932 2624 4959
rect 2658 4932 2697 4959
rect 2731 4932 2770 4959
rect 2804 4932 2843 4959
rect 2877 4932 2916 4959
rect 2950 4932 2989 4959
rect 3023 4932 3062 4959
rect 3096 4932 3135 4959
rect 3169 4932 3208 4959
rect 3242 4932 3281 4959
rect 3315 4932 3354 4959
rect 3388 4932 3427 4959
rect 3461 4932 3500 4959
rect 3534 4932 3573 4959
rect 3607 4932 3646 4959
rect 3680 4932 3719 4959
rect 3753 4932 3792 4959
rect 3826 4932 3865 4959
rect 3899 4932 3938 4959
rect 3972 4932 4011 4959
rect 4045 4932 4084 4959
rect 4118 4932 4157 4959
rect 4191 4932 4229 4959
rect 4263 4932 4301 4959
rect 4335 4932 4373 4959
rect 4407 4932 4445 4959
rect 4479 4932 4517 4959
rect 4551 4932 4589 4959
rect 4623 4932 4661 4959
rect 4695 4932 4733 4959
rect 4767 4932 4805 4959
rect 4839 4932 4877 4959
rect 4911 4932 4949 4959
rect 4983 4932 5021 4959
rect 5055 4932 5093 4959
rect 5127 4932 5165 4959
rect 5199 4932 5237 4959
rect 5271 4932 5309 4959
rect 5343 4932 5381 4959
rect 5415 4932 5453 4959
rect 5487 4932 5525 4959
rect 5559 4932 5597 4959
rect 5631 4932 5669 4959
rect 5703 4932 5741 4959
rect 5775 4932 5813 4959
rect 5847 4932 5885 4959
rect 5919 4932 5957 4959
rect 5991 4932 6029 4959
rect 6063 4932 6101 4959
rect 6135 4932 6173 4959
rect 6207 4932 6245 4959
rect 6279 4932 6317 4959
rect 6351 4932 6389 4959
rect 6423 4932 6461 4959
rect 6495 4932 6533 4959
rect 6567 4932 6605 4959
rect 6639 4932 6677 4959
rect 6711 4932 6749 4959
rect 6783 4932 6821 4959
rect 6855 4932 6893 4959
rect 6927 4932 6965 4959
rect 6999 4932 7037 4959
rect 7071 4932 7109 4959
rect 7143 4932 7181 4959
rect 7215 4932 7253 4959
rect 7287 4932 7325 4959
rect 7359 4932 7397 4959
rect 7431 4932 7469 4959
rect 7503 4932 7541 4959
rect 7575 4932 7613 4959
rect 7647 4932 7685 4959
rect 7719 4932 7757 4959
rect 7791 4932 7829 4959
rect 7863 4932 7901 4959
rect 7935 4932 7973 4959
rect 8007 4932 8045 4959
rect 8079 4932 8117 4959
rect 8151 4932 8189 4959
rect 8223 4932 8261 4959
rect 8295 4932 8333 4959
rect 8367 4932 8405 4959
rect 8439 4932 8477 4959
rect 8511 4932 8549 4959
rect 8583 4932 8621 4959
rect 8655 4932 8693 4959
rect 8727 4932 8765 4959
rect 8799 4932 8837 4959
rect 8871 4932 8909 4959
rect 8943 4932 8981 4959
rect 9015 4932 9053 4959
rect 9087 4932 9125 4959
rect 9159 4932 9197 4959
rect 9231 4932 9269 4959
rect 9303 4932 9341 4959
rect 9375 4932 9413 4959
rect 9447 4932 9485 4959
rect 9519 4932 9557 4959
rect 9591 4932 9629 4959
rect 9663 4932 9701 4959
rect 9735 4932 9773 4959
rect 9807 4932 9845 4959
rect 9879 4932 9917 4959
rect 9951 4932 9989 4959
rect 10023 4932 10061 4959
rect 10095 4932 10133 4959
rect 10167 4932 10205 4959
rect 10239 4932 10277 4959
rect 10311 4932 10349 4959
rect 10383 4932 10421 4959
rect 10455 4932 10493 4959
rect 10527 4932 10565 4959
rect 10599 4932 10637 4959
rect 10671 4932 10709 4959
rect 10743 4932 10781 4959
rect 10815 4932 10853 4959
rect 10887 4932 10925 4959
rect 10959 4932 10997 4959
rect 11031 4932 11069 4959
rect 11103 4932 11141 4959
rect 11175 4932 11213 4959
rect 11247 4932 11285 4959
rect 11319 4932 11357 4959
rect 11391 4932 11429 4959
rect 11463 4932 11501 4959
rect 11535 4932 11573 4959
rect 11607 4932 11645 4959
rect 11679 4932 11717 4959
rect 11751 4932 11789 4959
rect 11823 4932 11861 4959
rect 11895 4932 11933 4959
rect 11967 4932 12005 4959
rect 12039 4932 12077 4959
rect 12111 4932 12149 4959
rect 12183 4932 12221 4959
rect 12255 4932 12293 4959
rect 12327 4932 12365 4959
rect 12399 4932 12437 4959
rect 12471 4932 12509 4959
rect 12543 4932 12581 4959
rect 12615 4932 12653 4959
rect 12687 4932 12725 4959
rect 12759 4932 12797 4959
rect 12831 4932 12869 4959
rect 12903 4932 12941 4959
rect 12975 4932 13013 4959
rect 13047 4932 13085 4959
rect 13119 4932 13157 4959
rect 13191 4932 13229 4959
rect 13263 4932 13301 4959
rect 13335 4932 13373 4959
rect 13407 4932 13445 4959
rect 13479 4932 13517 4959
rect 13551 4932 13589 4959
rect 13623 4932 13661 4959
rect 13695 4932 13733 4959
rect 13767 4932 13805 4959
rect 13839 4932 13877 4959
rect 13911 4932 13949 4959
rect 13983 4932 14021 4959
rect 941 4898 979 4925
rect 1013 4925 1018 4932
rect 1085 4925 1091 4932
rect 1157 4925 1164 4932
rect 1229 4925 1237 4932
rect 1301 4925 1310 4932
rect 1373 4925 1383 4932
rect 1445 4925 1456 4932
rect 1517 4925 1529 4932
rect 1589 4925 1602 4932
rect 1661 4925 1675 4932
rect 1733 4925 1748 4932
rect 1805 4925 1821 4932
rect 1877 4925 1894 4932
rect 1949 4925 1967 4932
rect 2021 4925 2040 4932
rect 2093 4925 2113 4932
rect 2165 4925 2186 4932
rect 2237 4925 2259 4932
rect 2309 4925 2332 4932
rect 2381 4925 2405 4932
rect 2453 4925 2478 4932
rect 2525 4925 2551 4932
rect 2597 4925 2624 4932
rect 2669 4925 2697 4932
rect 2741 4925 2770 4932
rect 2813 4925 2843 4932
rect 2885 4925 2916 4932
rect 2957 4925 2989 4932
rect 3029 4925 3062 4932
rect 3101 4925 3135 4932
rect 3173 4925 3208 4932
rect 3245 4925 3281 4932
rect 3317 4925 3354 4932
rect 1013 4898 1051 4925
rect 1085 4898 1123 4925
rect 1157 4898 1195 4925
rect 1229 4898 1267 4925
rect 1301 4898 1339 4925
rect 1373 4898 1411 4925
rect 1445 4898 1483 4925
rect 1517 4898 1555 4925
rect 1589 4898 1627 4925
rect 1661 4898 1699 4925
rect 1733 4898 1771 4925
rect 1805 4898 1843 4925
rect 1877 4898 1915 4925
rect 1949 4898 1987 4925
rect 2021 4898 2059 4925
rect 2093 4898 2131 4925
rect 2165 4898 2203 4925
rect 2237 4898 2275 4925
rect 2309 4898 2347 4925
rect 2381 4898 2419 4925
rect 2453 4898 2491 4925
rect 2525 4898 2563 4925
rect 2597 4898 2635 4925
rect 2669 4898 2707 4925
rect 2741 4898 2779 4925
rect 2813 4898 2851 4925
rect 2885 4898 2923 4925
rect 2957 4898 2995 4925
rect 3029 4898 3067 4925
rect 3101 4898 3139 4925
rect 3173 4898 3211 4925
rect 3245 4898 3283 4925
rect 3317 4898 3355 4925
rect 3389 4898 3427 4932
rect 3461 4898 3499 4932
rect 3534 4925 3571 4932
rect 3607 4925 3643 4932
rect 3680 4925 3715 4932
rect 3753 4925 3787 4932
rect 3826 4925 3859 4932
rect 3899 4925 3931 4932
rect 3972 4925 4003 4932
rect 4045 4925 4075 4932
rect 4118 4925 4147 4932
rect 4191 4925 4219 4932
rect 4263 4925 4291 4932
rect 4335 4925 4363 4932
rect 4407 4925 4435 4932
rect 4479 4925 4507 4932
rect 4551 4925 4579 4932
rect 4623 4925 4651 4932
rect 4695 4925 4723 4932
rect 4767 4925 4795 4932
rect 4839 4925 4867 4932
rect 4911 4925 4939 4932
rect 4983 4925 5011 4932
rect 5055 4925 5083 4932
rect 5127 4925 5155 4932
rect 5199 4925 5227 4932
rect 5271 4925 5299 4932
rect 5343 4925 5371 4932
rect 5415 4925 5443 4932
rect 5487 4925 5515 4932
rect 5559 4925 5587 4932
rect 5631 4925 5659 4932
rect 5703 4925 5731 4932
rect 5775 4925 5803 4932
rect 5847 4925 5875 4932
rect 5919 4925 5947 4932
rect 5991 4925 6019 4932
rect 6063 4925 6091 4932
rect 6135 4925 6163 4932
rect 6207 4925 6235 4932
rect 6279 4925 6307 4932
rect 6351 4925 6379 4932
rect 6423 4925 6451 4932
rect 6495 4925 6523 4932
rect 6567 4925 6595 4932
rect 6639 4925 6667 4932
rect 6711 4925 6739 4932
rect 6783 4925 6811 4932
rect 6855 4925 6883 4932
rect 6927 4925 6955 4932
rect 6999 4925 7027 4932
rect 7071 4925 7099 4932
rect 7143 4925 7171 4932
rect 7215 4925 7243 4932
rect 7287 4925 7315 4932
rect 7359 4925 7387 4932
rect 7431 4925 7459 4932
rect 7503 4925 7531 4932
rect 7575 4925 7603 4932
rect 7647 4925 7675 4932
rect 7719 4925 7747 4932
rect 7791 4925 7819 4932
rect 7863 4925 7891 4932
rect 7935 4925 7963 4932
rect 8007 4925 8035 4932
rect 8079 4925 8107 4932
rect 8151 4925 8179 4932
rect 8223 4925 8251 4932
rect 8295 4925 8323 4932
rect 8367 4925 8395 4932
rect 8439 4925 8467 4932
rect 8511 4925 8539 4932
rect 8583 4925 8611 4932
rect 8655 4925 8683 4932
rect 8727 4925 8755 4932
rect 8799 4925 8827 4932
rect 8871 4925 8899 4932
rect 8943 4925 8971 4932
rect 9015 4925 9043 4932
rect 9087 4925 9115 4932
rect 9159 4925 9187 4932
rect 9231 4925 9259 4932
rect 9303 4925 9331 4932
rect 9375 4925 9403 4932
rect 9447 4925 9475 4932
rect 9519 4925 9547 4932
rect 9591 4925 9619 4932
rect 9663 4925 9691 4932
rect 9735 4925 9763 4932
rect 9807 4925 9835 4932
rect 9879 4925 9907 4932
rect 9951 4925 9979 4932
rect 10023 4925 10051 4932
rect 10095 4925 10123 4932
rect 10167 4925 10195 4932
rect 10239 4925 10267 4932
rect 10311 4925 10339 4932
rect 10383 4925 10411 4932
rect 10455 4925 10483 4932
rect 10527 4925 10555 4932
rect 10599 4925 10627 4932
rect 10671 4925 10699 4932
rect 10743 4925 10771 4932
rect 10815 4925 10843 4932
rect 10887 4925 10915 4932
rect 10959 4925 10987 4932
rect 11031 4925 11059 4932
rect 11103 4925 11131 4932
rect 11175 4925 11203 4932
rect 11247 4925 11275 4932
rect 11319 4925 11347 4932
rect 11391 4925 11419 4932
rect 11463 4925 11491 4932
rect 11535 4925 11563 4932
rect 11607 4925 11635 4932
rect 11679 4925 11707 4932
rect 11751 4925 11779 4932
rect 11823 4925 11851 4932
rect 11895 4925 11923 4932
rect 11967 4925 11995 4932
rect 12039 4925 12067 4932
rect 12111 4925 12139 4932
rect 12183 4925 12211 4932
rect 12255 4925 12283 4932
rect 12327 4925 12355 4932
rect 12399 4925 12427 4932
rect 12471 4925 12499 4932
rect 12543 4925 12571 4932
rect 12615 4925 12643 4932
rect 12687 4925 12715 4932
rect 12759 4925 12787 4932
rect 12831 4925 12859 4932
rect 12903 4925 12931 4932
rect 12975 4925 13003 4932
rect 13047 4925 13075 4932
rect 13119 4925 13147 4932
rect 13191 4925 13219 4932
rect 13263 4925 13291 4932
rect 13335 4925 13363 4932
rect 13407 4925 13436 4932
rect 13479 4925 13509 4932
rect 13551 4925 13582 4932
rect 13623 4925 13655 4932
rect 13695 4925 13728 4932
rect 13767 4925 13801 4932
rect 13839 4925 13874 4932
rect 13911 4925 13947 4932
rect 13983 4925 14020 4932
rect 14055 4925 14093 4959
rect 14127 4925 14165 4959
rect 14199 4932 14237 4959
rect 14271 4932 14309 4959
rect 14343 4932 14381 4959
rect 14415 4932 14453 4959
rect 14487 4932 14525 4959
rect 14559 4932 14597 4959
rect 14631 4932 14669 4959
rect 14703 4932 14741 4959
rect 14775 4958 14907 4959
rect 14775 4932 14832 4958
rect 14200 4925 14237 4932
rect 14273 4925 14309 4932
rect 14346 4925 14381 4932
rect 14419 4925 14453 4932
rect 14492 4925 14525 4932
rect 14565 4925 14597 4932
rect 14638 4925 14669 4932
rect 14711 4925 14741 4932
rect 3533 4898 3571 4925
rect 3605 4898 3643 4925
rect 3677 4898 3715 4925
rect 3749 4898 3787 4925
rect 3821 4898 3859 4925
rect 3893 4898 3931 4925
rect 3965 4898 4003 4925
rect 4037 4898 4075 4925
rect 4109 4898 4147 4925
rect 4181 4898 4219 4925
rect 4253 4898 4291 4925
rect 4325 4898 4363 4925
rect 4397 4898 4435 4925
rect 4469 4898 4507 4925
rect 4541 4898 4579 4925
rect 4613 4898 4651 4925
rect 4685 4898 4723 4925
rect 4757 4898 4795 4925
rect 4829 4898 4867 4925
rect 4901 4898 4939 4925
rect 4973 4898 5011 4925
rect 5045 4898 5083 4925
rect 5117 4898 5155 4925
rect 5189 4898 5227 4925
rect 5261 4898 5299 4925
rect 5333 4898 5371 4925
rect 5405 4898 5443 4925
rect 5477 4898 5515 4925
rect 5549 4898 5587 4925
rect 5621 4898 5659 4925
rect 5693 4898 5731 4925
rect 5765 4898 5803 4925
rect 5837 4898 5875 4925
rect 5909 4898 5947 4925
rect 5981 4898 6019 4925
rect 6053 4898 6091 4925
rect 6125 4898 6163 4925
rect 6197 4898 6235 4925
rect 6269 4898 6307 4925
rect 6341 4898 6379 4925
rect 6413 4898 6451 4925
rect 6485 4898 6523 4925
rect 6557 4898 6595 4925
rect 6629 4898 6667 4925
rect 6701 4898 6739 4925
rect 6773 4898 6811 4925
rect 6845 4898 6883 4925
rect 6917 4898 6955 4925
rect 6989 4898 7027 4925
rect 7061 4898 7099 4925
rect 7133 4898 7171 4925
rect 7205 4898 7243 4925
rect 7277 4898 7315 4925
rect 7349 4898 7387 4925
rect 7421 4898 7459 4925
rect 7493 4898 7531 4925
rect 7565 4898 7603 4925
rect 7637 4898 7675 4925
rect 7709 4898 7747 4925
rect 7781 4898 7819 4925
rect 7853 4898 7891 4925
rect 7925 4898 7963 4925
rect 7997 4898 8035 4925
rect 8069 4898 8107 4925
rect 8141 4898 8179 4925
rect 8213 4898 8251 4925
rect 8285 4898 8323 4925
rect 8357 4898 8395 4925
rect 8429 4898 8467 4925
rect 8501 4898 8539 4925
rect 8573 4898 8611 4925
rect 8645 4898 8683 4925
rect 8717 4898 8755 4925
rect 8789 4898 8827 4925
rect 8861 4898 8899 4925
rect 8933 4898 8971 4925
rect 9005 4898 9043 4925
rect 9077 4898 9115 4925
rect 9149 4898 9187 4925
rect 9221 4898 9259 4925
rect 9293 4898 9331 4925
rect 9365 4898 9403 4925
rect 9437 4898 9475 4925
rect 9509 4898 9547 4925
rect 9581 4898 9619 4925
rect 9653 4898 9691 4925
rect 9725 4898 9763 4925
rect 9797 4898 9835 4925
rect 9869 4898 9907 4925
rect 9941 4898 9979 4925
rect 10013 4898 10051 4925
rect 10085 4898 10123 4925
rect 10157 4898 10195 4925
rect 10229 4898 10267 4925
rect 10301 4898 10339 4925
rect 10373 4898 10411 4925
rect 10445 4898 10483 4925
rect 10517 4898 10555 4925
rect 10589 4898 10627 4925
rect 10661 4898 10699 4925
rect 10733 4898 10771 4925
rect 10805 4898 10843 4925
rect 10877 4898 10915 4925
rect 10949 4898 10987 4925
rect 11021 4898 11059 4925
rect 11093 4898 11131 4925
rect 11165 4898 11203 4925
rect 11237 4898 11275 4925
rect 11309 4898 11347 4925
rect 11381 4898 11419 4925
rect 11453 4898 11491 4925
rect 11525 4898 11563 4925
rect 11597 4898 11635 4925
rect 11669 4898 11707 4925
rect 11741 4898 11779 4925
rect 11813 4898 11851 4925
rect 11885 4898 11923 4925
rect 11957 4898 11995 4925
rect 12029 4898 12067 4925
rect 12101 4898 12139 4925
rect 12173 4898 12211 4925
rect 12245 4898 12283 4925
rect 12317 4898 12355 4925
rect 12389 4898 12427 4925
rect 12461 4898 12499 4925
rect 12533 4898 12571 4925
rect 12605 4898 12643 4925
rect 12677 4898 12715 4925
rect 12749 4898 12787 4925
rect 12821 4898 12859 4925
rect 12893 4898 12931 4925
rect 12965 4898 13003 4925
rect 13037 4898 13075 4925
rect 13109 4898 13147 4925
rect 13181 4898 13219 4925
rect 13253 4898 13291 4925
rect 13325 4898 13363 4925
rect 13397 4898 13436 4925
rect 13470 4898 13509 4925
rect 13543 4898 13582 4925
rect 13616 4898 13655 4925
rect 13689 4898 13728 4925
rect 13762 4898 13801 4925
rect 13835 4898 13874 4925
rect 13908 4898 13947 4925
rect 13981 4898 14020 4925
rect 14054 4898 14093 4925
rect 14127 4898 14166 4925
rect 14200 4898 14239 4925
rect 14273 4898 14312 4925
rect 14346 4898 14385 4925
rect 14419 4898 14458 4925
rect 14492 4898 14531 4925
rect 14565 4898 14604 4925
rect 14638 4898 14677 4925
rect 14711 4898 14750 4925
rect 14784 4898 14823 4932
rect 14866 4924 14907 4958
rect 14857 4898 14907 4924
rect 229 4886 14907 4898
rect 229 4883 14832 4886
rect 229 4859 269 4883
rect 229 4825 262 4859
rect 303 4849 329 4883
rect 296 4825 329 4849
rect 229 4810 329 4825
rect 229 4791 269 4810
rect 229 4757 262 4791
rect 303 4776 329 4810
rect 296 4757 329 4776
rect 229 4737 329 4757
rect 229 4723 269 4737
rect 229 4689 262 4723
rect 303 4703 329 4737
rect 296 4689 329 4703
rect 229 4664 329 4689
rect 229 4655 269 4664
rect 229 4621 262 4655
rect 303 4630 329 4664
rect 14807 4852 14832 4883
rect 14866 4859 14907 4886
rect 14807 4825 14840 4852
rect 14874 4825 14907 4859
rect 14807 4814 14907 4825
rect 14807 4780 14832 4814
rect 14866 4791 14907 4814
rect 14807 4757 14840 4780
rect 14874 4757 14907 4791
rect 14807 4742 14907 4757
rect 14807 4708 14832 4742
rect 14866 4723 14907 4742
rect 14807 4689 14840 4708
rect 14874 4689 14907 4723
rect 14807 4670 14907 4689
rect 296 4621 329 4630
rect 229 4591 329 4621
rect 229 4587 269 4591
rect 229 4553 262 4587
rect 303 4557 329 4591
rect 296 4553 329 4557
rect 229 4519 329 4553
rect 229 4485 262 4519
rect 296 4518 329 4519
rect 229 4484 269 4485
rect 303 4484 329 4518
rect 229 4451 329 4484
rect 229 4417 262 4451
rect 296 4445 329 4451
rect 229 4411 269 4417
rect 303 4411 329 4445
rect 229 4383 329 4411
rect 229 4349 262 4383
rect 296 4372 329 4383
rect 229 4338 269 4349
rect 303 4338 329 4372
rect 229 4315 329 4338
rect 229 4281 262 4315
rect 296 4299 329 4315
rect 229 4265 269 4281
rect 303 4265 329 4299
rect 229 4247 329 4265
rect 229 4213 262 4247
rect 296 4226 329 4247
rect 229 4192 269 4213
rect 303 4192 329 4226
rect 229 4179 329 4192
rect 229 4145 262 4179
rect 296 4153 329 4179
rect 229 4119 269 4145
rect 303 4119 329 4153
rect 229 4111 329 4119
rect 229 4077 262 4111
rect 296 4080 329 4111
rect 229 4046 269 4077
rect 303 4046 329 4080
rect 229 4043 329 4046
rect 229 4009 262 4043
rect 296 4009 329 4043
rect 229 4007 329 4009
rect 229 3975 269 4007
rect 229 3941 262 3975
rect 303 3973 329 4007
rect 296 3941 329 3973
rect 229 3934 329 3941
rect 229 3907 269 3934
rect 229 3873 262 3907
rect 303 3900 329 3934
rect 296 3873 329 3900
rect 229 3861 329 3873
rect 229 3839 269 3861
rect 229 3805 262 3839
rect 303 3827 329 3861
rect 296 3805 329 3827
rect 229 3788 329 3805
rect 229 3771 269 3788
rect 229 3737 262 3771
rect 303 3754 329 3788
rect 296 3737 329 3754
rect 229 3715 329 3737
rect 229 3703 269 3715
rect 229 3669 262 3703
rect 303 3681 329 3715
rect 296 3669 329 3681
rect 229 3642 329 3669
rect 229 3635 269 3642
rect 229 3601 262 3635
rect 303 3608 329 3642
rect 296 3601 329 3608
rect 229 3569 329 3601
rect 229 3567 269 3569
rect 229 3533 262 3567
rect 303 3535 329 3569
rect 296 3533 329 3535
rect 229 3499 329 3533
rect 229 3465 262 3499
rect 296 3496 329 3499
rect 229 3462 269 3465
rect 303 3462 329 3496
rect 229 3431 329 3462
rect 229 3397 262 3431
rect 296 3423 329 3431
rect 229 3389 269 3397
rect 303 3389 329 3423
rect 229 3363 329 3389
rect 229 3329 262 3363
rect 296 3350 329 3363
rect 229 3316 269 3329
rect 303 3316 329 3350
rect 229 3295 329 3316
rect 229 3261 262 3295
rect 296 3277 329 3295
rect 229 3243 269 3261
rect 303 3243 329 3277
rect 229 3227 329 3243
rect 229 3193 262 3227
rect 296 3204 329 3227
rect 229 3170 269 3193
rect 303 3170 329 3204
rect 229 3159 329 3170
rect 229 3125 262 3159
rect 296 3131 329 3159
rect 229 3097 269 3125
rect 303 3097 329 3131
rect 229 3091 329 3097
rect 229 3057 262 3091
rect 296 3058 329 3091
rect 229 3024 269 3057
rect 303 3024 329 3058
rect 229 3023 329 3024
rect 229 2989 262 3023
rect 296 2989 329 3023
rect 229 2985 329 2989
rect 229 2955 269 2985
rect 229 2921 262 2955
rect 303 2951 329 2985
rect 296 2921 329 2951
rect 229 2912 329 2921
rect 229 2887 269 2912
rect 229 2853 262 2887
rect 303 2878 329 2912
rect 296 2853 329 2878
rect 229 2839 329 2853
rect 229 2819 269 2839
rect 229 2785 262 2819
rect 303 2805 329 2839
rect 296 2785 329 2805
rect 229 2766 329 2785
rect 229 2751 269 2766
rect 229 2717 262 2751
rect 303 2732 329 2766
rect 296 2717 329 2732
rect 229 2693 329 2717
rect 229 2683 269 2693
rect 229 2649 262 2683
rect 303 2659 329 2693
rect 296 2649 329 2659
rect 229 2620 329 2649
rect 229 2615 269 2620
rect 229 2581 262 2615
rect 303 2586 329 2620
rect 296 2581 329 2586
rect 229 2547 329 2581
rect 229 2513 262 2547
rect 303 2513 329 2547
rect 229 2479 329 2513
rect 229 2445 262 2479
rect 296 2474 329 2479
rect 229 2440 269 2445
rect 303 2440 329 2474
rect 229 2411 329 2440
rect 229 2377 262 2411
rect 296 2401 329 2411
rect 229 2367 269 2377
rect 303 2367 329 2401
rect 229 2343 329 2367
rect 229 2309 262 2343
rect 296 2328 329 2343
rect 229 2294 269 2309
rect 303 2294 329 2328
rect 229 2275 329 2294
rect 229 2241 262 2275
rect 296 2255 329 2275
rect 229 2221 269 2241
rect 303 2221 329 2255
rect 229 2207 329 2221
rect 229 2173 262 2207
rect 296 2182 329 2207
rect 229 2148 269 2173
rect 303 2148 329 2182
rect 229 2139 329 2148
rect 229 2105 262 2139
rect 296 2109 329 2139
rect 229 2075 269 2105
rect 303 2075 329 2109
rect 229 2071 329 2075
rect 229 2037 262 2071
rect 296 2037 329 2071
rect 229 2036 329 2037
rect 229 2003 269 2036
rect 229 1969 262 2003
rect 303 2002 329 2036
rect 296 1969 329 2002
rect 229 1963 329 1969
rect 229 1935 269 1963
rect 229 1901 262 1935
rect 303 1929 329 1963
rect 296 1901 329 1929
rect 229 1890 329 1901
rect 229 1867 269 1890
rect 229 1833 262 1867
rect 303 1856 329 1890
rect 296 1833 329 1856
rect 229 1817 329 1833
rect 229 1799 269 1817
rect 229 1765 262 1799
rect 303 1783 329 1817
rect 296 1765 329 1783
rect 229 1744 329 1765
rect 229 1731 269 1744
rect 229 1697 262 1731
rect 303 1710 329 1744
rect 296 1697 329 1710
rect 229 1671 329 1697
rect 229 1663 269 1671
rect 229 1629 262 1663
rect 303 1637 329 1671
rect 296 1629 329 1637
rect 229 1598 329 1629
rect 229 1595 269 1598
rect 229 1561 262 1595
rect 303 1564 329 1598
rect 296 1561 329 1564
rect 229 1527 329 1561
rect 229 1493 262 1527
rect 296 1525 329 1527
rect 229 1491 269 1493
rect 303 1491 329 1525
rect 229 1459 329 1491
rect 229 1425 262 1459
rect 296 1452 329 1459
rect 229 1418 269 1425
rect 303 1418 329 1452
rect 229 1391 329 1418
rect 229 1357 262 1391
rect 296 1379 329 1391
rect 229 1345 269 1357
rect 303 1345 329 1379
rect 229 1323 329 1345
rect 229 1289 262 1323
rect 296 1306 329 1323
rect 229 1272 269 1289
rect 303 1272 329 1306
rect 229 1255 329 1272
rect 229 1221 262 1255
rect 296 1233 329 1255
rect 229 1199 269 1221
rect 303 1199 329 1233
rect 229 1187 329 1199
rect 229 1153 262 1187
rect 296 1159 329 1187
rect 229 1125 269 1153
rect 303 1125 329 1159
rect 229 1119 329 1125
rect 229 1085 262 1119
rect 296 1085 329 1119
rect 229 1051 269 1085
rect 303 1051 329 1085
rect 229 1017 262 1051
rect 296 1017 329 1051
rect 229 1011 329 1017
rect 229 983 269 1011
rect 229 949 262 983
rect 303 977 329 1011
rect 296 949 329 977
rect 229 937 329 949
rect 229 915 269 937
rect 229 881 262 915
rect 303 903 329 937
rect 296 881 329 903
rect 229 863 329 881
rect 229 847 269 863
rect 229 813 262 847
rect 303 829 329 863
rect 296 813 329 829
rect 229 789 329 813
rect 229 779 269 789
rect 229 745 262 779
rect 303 755 329 789
rect 296 745 329 755
rect 229 715 329 745
rect 229 711 269 715
rect 229 677 262 711
rect 303 681 329 715
rect 296 677 329 681
rect 229 643 329 677
rect 482 4638 14653 4653
rect 482 4619 584 4638
rect 482 4585 497 4619
rect 531 4585 584 4619
rect 10410 4606 10445 4638
rect 10479 4606 10514 4638
rect 10548 4606 10583 4638
rect 10617 4606 10652 4638
rect 10686 4606 10721 4638
rect 10755 4606 10790 4638
rect 10824 4606 10859 4638
rect 10893 4606 10928 4638
rect 10962 4606 10997 4638
rect 11031 4606 11066 4638
rect 11100 4606 11135 4638
rect 11169 4606 11204 4638
rect 11238 4606 11273 4638
rect 11307 4606 11342 4638
rect 11376 4606 11411 4638
rect 11445 4606 11480 4638
rect 11514 4606 11549 4638
rect 11583 4606 11618 4638
rect 11652 4606 11687 4638
rect 11721 4606 11756 4638
rect 11790 4606 11825 4638
rect 11859 4606 11894 4638
rect 11928 4606 11963 4638
rect 11997 4606 12032 4638
rect 12066 4606 12101 4638
rect 12135 4606 12170 4638
rect 12204 4606 12239 4638
rect 12273 4606 12308 4638
rect 12342 4606 12377 4638
rect 12411 4606 12446 4638
rect 12480 4606 12515 4638
rect 12549 4606 12584 4638
rect 12618 4606 12653 4638
rect 12687 4606 12722 4638
rect 12756 4606 12791 4638
rect 12825 4606 12860 4638
rect 12894 4606 12929 4638
rect 12963 4606 12998 4638
rect 13032 4606 13067 4638
rect 13101 4606 13136 4638
rect 13170 4606 13205 4638
rect 13239 4606 13274 4638
rect 13308 4606 13343 4638
rect 13377 4606 13412 4638
rect 13446 4606 13481 4638
rect 13515 4606 13550 4638
rect 13584 4606 13619 4638
rect 13653 4606 13688 4638
rect 13722 4606 13757 4638
rect 13791 4606 13826 4638
rect 13860 4606 13895 4638
rect 13929 4606 13964 4638
rect 13998 4606 14033 4638
rect 14067 4606 14102 4638
rect 14136 4606 14171 4638
rect 14205 4606 14240 4638
rect 14274 4606 14309 4638
rect 14343 4606 14378 4638
rect 14412 4606 14447 4638
rect 482 4570 584 4585
rect 14207 4604 14240 4606
rect 14280 4604 14309 4606
rect 14353 4604 14378 4606
rect 14426 4604 14447 4606
rect 14481 4604 14516 4638
rect 14550 4604 14585 4638
rect 14619 4604 14653 4638
rect 14207 4572 14246 4604
rect 14280 4572 14319 4604
rect 14353 4572 14392 4604
rect 14426 4572 14653 4604
rect 14207 4570 14653 4572
rect 482 4549 565 4570
rect 482 4515 497 4549
rect 531 4536 565 4549
rect 531 4515 633 4536
rect 482 4498 633 4515
rect 14225 4536 14260 4570
rect 14294 4536 14329 4570
rect 14363 4536 14398 4570
rect 14432 4536 14467 4570
rect 14501 4536 14536 4570
rect 14570 4551 14653 4570
rect 14207 4534 14536 4536
rect 14207 4502 14246 4534
rect 14280 4502 14319 4534
rect 14353 4502 14392 4534
rect 14426 4502 14536 4534
rect 14226 4500 14246 4502
rect 14295 4500 14319 4502
rect 14364 4500 14392 4502
rect 482 4479 565 4498
rect 482 4445 497 4479
rect 531 4464 565 4479
rect 599 4468 633 4498
rect 12363 4468 12398 4500
rect 12432 4468 12467 4500
rect 12501 4468 12536 4500
rect 12570 4468 12605 4500
rect 12639 4468 12674 4500
rect 12708 4468 12743 4500
rect 12777 4468 12812 4500
rect 12846 4468 12881 4500
rect 12915 4468 12950 4500
rect 12984 4468 13019 4500
rect 13053 4468 13088 4500
rect 13122 4468 13157 4500
rect 13191 4468 13226 4500
rect 13260 4468 13295 4500
rect 13329 4468 13364 4500
rect 13398 4468 13433 4500
rect 13467 4468 13502 4500
rect 13536 4468 13571 4500
rect 13605 4468 13640 4500
rect 13674 4468 13709 4500
rect 13743 4468 13778 4500
rect 13812 4468 13847 4500
rect 13881 4468 13916 4500
rect 13950 4468 13985 4500
rect 14019 4468 14054 4500
rect 14088 4468 14123 4500
rect 14157 4468 14192 4500
rect 14226 4468 14261 4500
rect 14295 4468 14330 4500
rect 14364 4468 14399 4500
rect 14433 4468 14468 4502
rect 599 4464 14468 4468
rect 531 4456 14468 4464
rect 531 4445 674 4456
rect 708 4453 14428 4456
rect 708 4445 780 4453
rect 482 4429 674 4445
rect 482 4426 633 4429
rect 482 4409 529 4426
rect 482 4375 497 4409
rect 563 4392 565 4426
rect 599 4392 601 4426
rect 667 4395 674 4429
rect 635 4392 674 4395
rect 531 4375 674 4392
rect 482 4356 674 4375
rect 482 4354 633 4356
rect 482 4351 565 4354
rect 482 4339 529 4351
rect 482 4305 497 4339
rect 563 4320 565 4351
rect 599 4351 633 4354
rect 599 4320 601 4351
rect 667 4322 674 4356
rect 563 4317 601 4320
rect 635 4317 674 4322
rect 531 4305 674 4317
rect 482 4283 674 4305
rect 482 4282 633 4283
rect 482 4276 565 4282
rect 482 4269 529 4276
rect 482 4235 497 4269
rect 563 4248 565 4276
rect 599 4276 633 4282
rect 599 4248 601 4276
rect 667 4249 674 4283
rect 563 4242 601 4248
rect 635 4242 674 4249
rect 531 4235 674 4242
rect 482 4211 674 4235
rect 482 4210 633 4211
rect 482 4201 565 4210
rect 482 4199 529 4201
rect 482 4165 497 4199
rect 563 4176 565 4201
rect 599 4201 633 4210
rect 599 4176 601 4201
rect 667 4177 674 4211
rect 563 4167 601 4176
rect 635 4167 674 4177
rect 531 4165 674 4167
rect 482 4139 674 4165
rect 482 4138 633 4139
rect 482 4129 565 4138
rect 482 4095 497 4129
rect 531 4126 565 4129
rect 563 4104 565 4126
rect 599 4126 633 4138
rect 599 4104 601 4126
rect 667 4105 674 4139
rect 482 4092 529 4095
rect 563 4092 601 4104
rect 635 4092 674 4105
rect 482 4067 674 4092
rect 14356 4432 14428 4453
rect 14390 4398 14428 4432
rect 14462 4426 14468 4456
rect 14356 4359 14428 4398
rect 14390 4325 14428 4359
rect 482 4066 633 4067
rect 482 4059 565 4066
rect 482 4025 497 4059
rect 531 4052 565 4059
rect 563 4032 565 4052
rect 599 4052 633 4066
rect 599 4032 601 4052
rect 667 4033 674 4067
rect 482 4018 529 4025
rect 563 4018 601 4032
rect 635 4018 674 4033
rect 482 3995 674 4018
rect 482 3994 633 3995
rect 482 3989 565 3994
rect 482 3955 497 3989
rect 531 3978 565 3989
rect 563 3960 565 3978
rect 599 3978 633 3994
rect 599 3960 601 3978
rect 667 3961 674 3995
rect 482 3944 529 3955
rect 563 3944 601 3960
rect 635 3944 674 3961
rect 482 3923 674 3944
rect 482 3922 633 3923
rect 482 3920 565 3922
rect 482 3886 497 3920
rect 531 3904 565 3920
rect 563 3888 565 3904
rect 599 3904 633 3922
rect 599 3888 601 3904
rect 667 3889 674 3923
rect 482 3870 529 3886
rect 563 3870 601 3888
rect 635 3870 674 3889
rect 482 3851 674 3870
rect 482 3817 497 3851
rect 531 3817 565 3851
rect 599 3817 633 3851
rect 667 3817 674 3851
rect 482 3794 674 3817
rect 482 3760 529 3794
rect 563 3760 601 3794
rect 635 3760 674 3794
rect 482 3749 674 3760
rect 482 3715 497 3749
rect 531 3720 565 3749
rect 563 3715 565 3720
rect 599 3720 633 3749
rect 599 3715 601 3720
rect 667 3715 674 3749
rect 482 3686 529 3715
rect 563 3686 601 3715
rect 635 3686 674 3715
rect 482 3680 674 3686
rect 482 3646 497 3680
rect 531 3646 565 3680
rect 599 3646 633 3680
rect 667 3646 674 3680
rect 482 3612 529 3646
rect 563 3612 601 3646
rect 635 3612 674 3646
rect 482 3611 674 3612
rect 482 3577 497 3611
rect 531 3577 565 3611
rect 599 3577 633 3611
rect 667 3577 674 3611
rect 482 3572 674 3577
rect 482 3542 529 3572
rect 563 3542 601 3572
rect 635 3542 674 3572
rect 482 3508 497 3542
rect 563 3538 565 3542
rect 531 3508 565 3538
rect 599 3538 601 3542
rect 599 3508 633 3538
rect 667 3508 674 3542
rect 482 3498 674 3508
rect 482 3473 529 3498
rect 563 3473 601 3498
rect 635 3473 674 3498
rect 482 3439 497 3473
rect 563 3464 565 3473
rect 531 3439 565 3464
rect 599 3464 601 3473
rect 599 3439 633 3464
rect 667 3439 674 3473
rect 482 3424 674 3439
rect 482 3404 529 3424
rect 563 3404 601 3424
rect 635 3404 674 3424
rect 482 3370 497 3404
rect 563 3390 565 3404
rect 531 3370 565 3390
rect 599 3390 601 3404
rect 599 3370 633 3390
rect 667 3370 674 3404
rect 482 3350 674 3370
rect 482 3335 529 3350
rect 563 3335 601 3350
rect 635 3335 674 3350
rect 482 3301 497 3335
rect 563 3316 565 3335
rect 531 3301 565 3316
rect 599 3316 601 3335
rect 599 3301 633 3316
rect 667 3301 674 3335
rect 482 3276 674 3301
rect 482 3266 529 3276
rect 563 3266 601 3276
rect 635 3266 674 3276
rect 482 3232 497 3266
rect 563 3242 565 3266
rect 531 3232 565 3242
rect 599 3242 601 3266
rect 599 3232 633 3242
rect 667 3232 674 3266
rect 482 3202 674 3232
rect 482 3197 529 3202
rect 563 3197 601 3202
rect 635 3197 674 3202
rect 482 3163 497 3197
rect 563 3168 565 3197
rect 531 3163 565 3168
rect 599 3168 601 3197
rect 599 3163 633 3168
rect 667 3163 674 3197
rect 482 3128 674 3163
rect 482 3094 497 3128
rect 563 3094 565 3128
rect 599 3094 601 3128
rect 667 3094 674 3128
rect 482 3059 674 3094
rect 482 3025 497 3059
rect 531 3054 565 3059
rect 563 3025 565 3054
rect 599 3054 633 3059
rect 599 3025 601 3054
rect 667 3025 674 3059
rect 482 3020 529 3025
rect 563 3020 601 3025
rect 635 3020 674 3025
rect 482 2990 674 3020
rect 482 2956 497 2990
rect 531 2980 565 2990
rect 563 2956 565 2980
rect 599 2980 633 2990
rect 599 2956 601 2980
rect 667 2956 674 2990
rect 482 2946 529 2956
rect 563 2946 601 2956
rect 635 2946 674 2956
rect 482 2921 674 2946
rect 482 2887 497 2921
rect 531 2906 565 2921
rect 563 2887 565 2906
rect 599 2906 633 2921
rect 599 2887 601 2906
rect 667 2887 674 2921
rect 482 2872 529 2887
rect 563 2872 601 2887
rect 635 2872 674 2887
rect 482 2852 674 2872
rect 482 2818 497 2852
rect 531 2832 565 2852
rect 563 2818 565 2832
rect 599 2832 633 2852
rect 599 2818 601 2832
rect 667 2818 674 2852
rect 482 2798 529 2818
rect 563 2798 601 2818
rect 635 2798 674 2818
rect 482 2783 674 2798
rect 482 2749 497 2783
rect 531 2758 565 2783
rect 563 2749 565 2758
rect 599 2758 633 2783
rect 599 2749 601 2758
rect 667 2749 674 2783
rect 482 2724 529 2749
rect 563 2724 601 2749
rect 635 2724 674 2749
rect 482 2714 674 2724
rect 482 2680 497 2714
rect 531 2684 565 2714
rect 563 2680 565 2684
rect 599 2684 633 2714
rect 599 2680 601 2684
rect 667 2680 674 2714
rect 482 2650 529 2680
rect 563 2650 601 2680
rect 635 2650 674 2680
rect 482 2645 674 2650
rect 482 2611 497 2645
rect 531 2611 565 2645
rect 599 2611 633 2645
rect 667 2611 674 2645
rect 482 2610 674 2611
rect 482 2576 529 2610
rect 563 2576 601 2610
rect 635 2576 674 2610
rect 482 2542 497 2576
rect 531 2542 565 2576
rect 599 2542 633 2576
rect 667 2542 674 2576
rect 482 2536 674 2542
rect 482 2507 529 2536
rect 563 2507 601 2536
rect 635 2507 674 2536
rect 482 2473 497 2507
rect 563 2502 565 2507
rect 531 2473 565 2502
rect 599 2502 601 2507
rect 599 2473 633 2502
rect 667 2473 674 2507
rect 482 2462 674 2473
rect 482 2438 529 2462
rect 563 2438 601 2462
rect 635 2438 674 2462
rect 482 2404 497 2438
rect 563 2428 565 2438
rect 531 2404 565 2428
rect 599 2428 601 2438
rect 599 2404 633 2428
rect 667 2404 674 2438
rect 482 2389 674 2404
rect 482 2369 529 2389
rect 563 2369 601 2389
rect 635 2369 674 2389
rect 482 2335 497 2369
rect 563 2355 565 2369
rect 531 2335 565 2355
rect 599 2355 601 2369
rect 599 2335 633 2355
rect 667 2335 674 2369
rect 482 2316 674 2335
rect 482 2300 529 2316
rect 563 2300 601 2316
rect 635 2300 674 2316
rect 482 2266 497 2300
rect 563 2282 565 2300
rect 531 2266 565 2282
rect 599 2282 601 2300
rect 599 2266 633 2282
rect 667 2266 674 2300
rect 482 2243 674 2266
rect 482 2231 529 2243
rect 563 2231 601 2243
rect 635 2231 674 2243
rect 482 2197 497 2231
rect 563 2209 565 2231
rect 531 2197 565 2209
rect 599 2209 601 2231
rect 599 2197 633 2209
rect 667 2197 674 2231
rect 482 2170 674 2197
rect 482 2163 529 2170
rect 482 2129 497 2163
rect 563 2162 601 2170
rect 635 2162 674 2170
rect 563 2136 565 2162
rect 531 2129 565 2136
rect 482 2128 565 2129
rect 599 2136 601 2162
rect 599 2128 633 2136
rect 667 2128 674 2162
rect 482 2097 674 2128
rect 482 2095 529 2097
rect 482 2061 497 2095
rect 563 2093 601 2097
rect 635 2093 674 2097
rect 563 2063 565 2093
rect 531 2061 565 2063
rect 482 2059 565 2061
rect 599 2063 601 2093
rect 599 2059 633 2063
rect 667 2059 674 2093
rect 482 2027 674 2059
rect 482 1993 497 2027
rect 531 2024 674 2027
rect 482 1990 529 1993
rect 563 1990 565 2024
rect 599 1990 601 2024
rect 667 1990 674 2024
rect 482 1959 674 1990
rect 482 1925 497 1959
rect 531 1955 674 1959
rect 531 1951 565 1955
rect 482 1917 529 1925
rect 563 1921 565 1951
rect 599 1951 633 1955
rect 599 1921 601 1951
rect 667 1921 674 1955
rect 563 1917 601 1921
rect 635 1917 674 1921
rect 482 1891 674 1917
rect 482 1857 497 1891
rect 531 1886 674 1891
rect 531 1878 565 1886
rect 482 1844 529 1857
rect 563 1852 565 1878
rect 599 1878 633 1886
rect 599 1852 601 1878
rect 667 1852 674 1886
rect 563 1844 601 1852
rect 635 1844 674 1852
rect 482 1823 674 1844
rect 482 1789 497 1823
rect 531 1817 674 1823
rect 531 1805 565 1817
rect 482 1771 529 1789
rect 563 1783 565 1805
rect 599 1805 633 1817
rect 599 1783 601 1805
rect 667 1783 674 1817
rect 563 1771 601 1783
rect 635 1771 674 1783
rect 482 1755 674 1771
rect 482 1721 497 1755
rect 531 1748 674 1755
rect 531 1732 565 1748
rect 482 1698 529 1721
rect 563 1714 565 1732
rect 599 1732 633 1748
rect 599 1714 601 1732
rect 667 1714 674 1748
rect 563 1698 601 1714
rect 635 1698 674 1714
rect 482 1687 674 1698
rect 482 1653 497 1687
rect 531 1679 674 1687
rect 531 1659 565 1679
rect 482 1625 529 1653
rect 563 1645 565 1659
rect 599 1659 633 1679
rect 599 1645 601 1659
rect 667 1645 674 1679
rect 563 1625 601 1645
rect 635 1625 674 1645
rect 482 1619 674 1625
rect 482 1585 497 1619
rect 531 1610 674 1619
rect 531 1586 565 1610
rect 482 1552 529 1585
rect 563 1576 565 1586
rect 599 1586 633 1610
rect 599 1576 601 1586
rect 667 1576 674 1610
rect 563 1552 601 1576
rect 635 1552 674 1576
rect 482 1551 674 1552
rect 482 1517 497 1551
rect 531 1541 674 1551
rect 531 1517 565 1541
rect 482 1513 565 1517
rect 482 1483 529 1513
rect 563 1507 565 1513
rect 599 1513 633 1541
rect 599 1507 601 1513
rect 667 1507 674 1541
rect 482 1449 497 1483
rect 563 1479 601 1507
rect 635 1479 674 1507
rect 531 1472 674 1479
rect 531 1449 565 1472
rect 482 1440 565 1449
rect 482 1415 529 1440
rect 563 1438 565 1440
rect 599 1440 633 1472
rect 599 1438 601 1440
rect 667 1438 674 1472
rect 482 1381 497 1415
rect 563 1406 601 1438
rect 635 1406 674 1438
rect 531 1403 674 1406
rect 531 1381 565 1403
rect 482 1369 565 1381
rect 599 1369 633 1403
rect 667 1369 674 1403
rect 482 1367 674 1369
rect 482 1347 529 1367
rect 482 1313 497 1347
rect 563 1334 601 1367
rect 635 1334 674 1367
rect 563 1333 565 1334
rect 531 1313 565 1333
rect 482 1300 565 1313
rect 599 1333 601 1334
rect 599 1300 633 1333
rect 667 1300 674 1334
rect 482 1294 674 1300
rect 482 1279 529 1294
rect 482 1245 497 1279
rect 563 1265 601 1294
rect 635 1265 674 1294
rect 563 1260 565 1265
rect 531 1245 565 1260
rect 482 1231 565 1245
rect 599 1260 601 1265
rect 599 1231 633 1260
rect 667 1231 674 1265
rect 482 1221 674 1231
rect 482 1211 529 1221
rect 482 1177 497 1211
rect 563 1196 601 1221
rect 635 1196 674 1221
rect 563 1187 565 1196
rect 531 1177 565 1187
rect 482 1162 565 1177
rect 599 1187 601 1196
rect 599 1162 633 1187
rect 667 1162 674 1196
rect 482 1148 674 1162
rect 482 1143 529 1148
rect 482 1109 497 1143
rect 563 1127 601 1148
rect 635 1127 674 1148
rect 563 1114 565 1127
rect 531 1109 565 1114
rect 482 1093 565 1109
rect 599 1114 601 1127
rect 599 1093 633 1114
rect 667 1093 674 1127
rect 482 1075 674 1093
rect 482 1041 497 1075
rect 563 1058 601 1075
rect 635 1058 674 1075
rect 563 1041 565 1058
rect 482 1024 565 1041
rect 599 1041 601 1058
rect 599 1024 633 1041
rect 667 1024 674 1058
rect 482 1007 674 1024
rect 482 973 497 1007
rect 531 1002 674 1007
rect 563 989 601 1002
rect 635 989 674 1002
rect 482 968 529 973
rect 563 968 565 989
rect 482 955 565 968
rect 599 968 601 989
rect 599 955 633 968
rect 667 955 674 989
rect 482 939 674 955
rect 482 769 497 939
rect 531 929 674 939
rect 563 920 601 929
rect 635 920 674 929
rect 667 894 674 920
rect 881 4308 1001 4324
rect 881 4274 924 4308
rect 958 4274 1001 4308
rect 881 4234 1001 4274
rect 881 4200 924 4234
rect 958 4200 1001 4234
rect 881 3104 1001 4200
rect 1311 4308 1431 4324
rect 1311 4274 1354 4308
rect 1388 4274 1431 4308
rect 1311 4234 1431 4274
rect 1311 4200 1354 4234
rect 1388 4200 1431 4234
rect 881 3070 924 3104
rect 958 3070 1001 3104
rect 881 3026 1001 3070
rect 881 2992 924 3026
rect 958 2992 1001 3026
rect 881 2948 1001 2992
rect 881 2914 924 2948
rect 958 2914 1001 2948
rect 881 2870 1001 2914
rect 881 2836 924 2870
rect 958 2836 1001 2870
rect 881 2792 1001 2836
rect 881 2758 924 2792
rect 958 2758 1001 2792
rect 881 2713 1001 2758
rect 881 2679 924 2713
rect 958 2679 1001 2713
rect 881 2634 1001 2679
rect 881 2600 924 2634
rect 958 2600 1001 2634
rect 881 1504 1001 2600
rect 1066 4064 1067 4098
rect 1101 4082 1139 4098
rect 1101 4064 1103 4082
rect 1066 4048 1103 4064
rect 1137 4064 1139 4082
rect 1173 4082 1211 4098
rect 1173 4064 1175 4082
rect 1137 4048 1175 4064
rect 1209 4064 1211 4082
rect 1245 4064 1246 4098
rect 1209 4048 1246 4064
rect 1066 4025 1246 4048
rect 1066 3991 1067 4025
rect 1101 4014 1139 4025
rect 1101 3991 1103 4014
rect 1066 3980 1103 3991
rect 1137 3991 1139 4014
rect 1173 4014 1211 4025
rect 1173 3991 1175 4014
rect 1137 3980 1175 3991
rect 1209 3991 1211 4014
rect 1245 3991 1246 4025
rect 1209 3980 1246 3991
rect 1066 3952 1246 3980
rect 1066 3918 1067 3952
rect 1101 3946 1139 3952
rect 1101 3918 1103 3946
rect 1066 3912 1103 3918
rect 1137 3918 1139 3946
rect 1173 3946 1211 3952
rect 1173 3918 1175 3946
rect 1137 3912 1175 3918
rect 1209 3918 1211 3946
rect 1245 3918 1246 3952
rect 1209 3912 1246 3918
rect 1066 3879 1246 3912
rect 1066 3845 1067 3879
rect 1101 3878 1139 3879
rect 1101 3845 1103 3878
rect 1066 3844 1103 3845
rect 1137 3845 1139 3878
rect 1173 3878 1211 3879
rect 1173 3845 1175 3878
rect 1137 3844 1175 3845
rect 1209 3845 1211 3878
rect 1245 3845 1246 3879
rect 1209 3844 1246 3845
rect 1066 3810 1246 3844
rect 1066 3806 1103 3810
rect 1066 3772 1067 3806
rect 1101 3776 1103 3806
rect 1137 3806 1175 3810
rect 1137 3776 1139 3806
rect 1101 3772 1139 3776
rect 1173 3776 1175 3806
rect 1209 3806 1246 3810
rect 1209 3776 1211 3806
rect 1173 3772 1211 3776
rect 1245 3772 1246 3806
rect 1066 3742 1246 3772
rect 1066 3733 1103 3742
rect 1066 3699 1067 3733
rect 1101 3708 1103 3733
rect 1137 3733 1175 3742
rect 1137 3708 1139 3733
rect 1101 3699 1139 3708
rect 1173 3708 1175 3733
rect 1209 3733 1246 3742
rect 1209 3708 1211 3733
rect 1173 3699 1211 3708
rect 1245 3699 1246 3733
rect 1066 3674 1246 3699
rect 1066 3660 1103 3674
rect 1066 3626 1067 3660
rect 1101 3640 1103 3660
rect 1137 3660 1175 3674
rect 1137 3640 1139 3660
rect 1101 3626 1139 3640
rect 1173 3640 1175 3660
rect 1209 3660 1246 3674
rect 1209 3640 1211 3660
rect 1173 3626 1211 3640
rect 1245 3626 1246 3660
rect 1066 3606 1246 3626
rect 1066 3587 1103 3606
rect 1066 3553 1067 3587
rect 1101 3572 1103 3587
rect 1137 3587 1175 3606
rect 1137 3572 1139 3587
rect 1101 3553 1139 3572
rect 1173 3572 1175 3587
rect 1209 3587 1246 3606
rect 1209 3572 1211 3587
rect 1173 3553 1211 3572
rect 1245 3553 1246 3587
rect 1066 3538 1246 3553
rect 1066 3514 1103 3538
rect 1066 3480 1067 3514
rect 1101 3504 1103 3514
rect 1137 3514 1175 3538
rect 1137 3504 1139 3514
rect 1101 3480 1139 3504
rect 1173 3504 1175 3514
rect 1209 3514 1246 3538
rect 1209 3504 1211 3514
rect 1173 3480 1211 3504
rect 1245 3480 1246 3514
rect 1066 3470 1246 3480
rect 1066 3441 1103 3470
rect 1066 3407 1067 3441
rect 1101 3436 1103 3441
rect 1137 3441 1175 3470
rect 1137 3436 1139 3441
rect 1101 3407 1139 3436
rect 1173 3436 1175 3441
rect 1209 3441 1246 3470
rect 1209 3436 1211 3441
rect 1173 3407 1211 3436
rect 1245 3407 1246 3441
rect 1066 3402 1246 3407
rect 1066 3368 1103 3402
rect 1137 3368 1175 3402
rect 1209 3368 1246 3402
rect 1066 3334 1067 3368
rect 1101 3334 1139 3368
rect 1173 3334 1211 3368
rect 1245 3334 1246 3368
rect 1066 3300 1103 3334
rect 1137 3300 1175 3334
rect 1209 3300 1246 3334
rect 1066 3295 1246 3300
rect 1066 3261 1067 3295
rect 1101 3266 1139 3295
rect 1101 3261 1103 3266
rect 1066 3232 1103 3261
rect 1137 3261 1139 3266
rect 1173 3266 1211 3295
rect 1173 3261 1175 3266
rect 1137 3232 1175 3261
rect 1209 3261 1211 3266
rect 1245 3261 1246 3295
rect 1209 3232 1246 3261
rect 1066 3222 1246 3232
rect 1066 3188 1067 3222
rect 1101 3198 1139 3222
rect 1101 3188 1103 3198
rect 1066 3164 1103 3188
rect 1137 3188 1139 3198
rect 1173 3198 1211 3222
rect 1173 3188 1175 3198
rect 1137 3164 1175 3188
rect 1209 3188 1211 3198
rect 1245 3188 1246 3222
rect 1209 3164 1246 3188
rect 1066 3149 1246 3164
rect 1066 3115 1067 3149
rect 1101 3115 1139 3149
rect 1173 3115 1211 3149
rect 1245 3115 1246 3149
rect 1066 3076 1246 3115
rect 1066 3042 1067 3076
rect 1101 3042 1139 3076
rect 1173 3042 1211 3076
rect 1245 3042 1246 3076
rect 1066 3003 1246 3042
rect 1066 2969 1067 3003
rect 1101 2969 1139 3003
rect 1173 2969 1211 3003
rect 1245 2969 1246 3003
rect 1066 2930 1246 2969
rect 1066 2896 1067 2930
rect 1101 2896 1139 2930
rect 1173 2896 1211 2930
rect 1245 2896 1246 2930
rect 1066 2857 1246 2896
rect 1066 2823 1067 2857
rect 1101 2823 1139 2857
rect 1173 2823 1211 2857
rect 1245 2823 1246 2857
rect 1066 2784 1246 2823
rect 1066 2750 1067 2784
rect 1101 2750 1139 2784
rect 1173 2750 1211 2784
rect 1245 2750 1246 2784
rect 1066 2711 1246 2750
rect 1066 2677 1067 2711
rect 1101 2677 1139 2711
rect 1173 2677 1211 2711
rect 1245 2677 1246 2711
rect 1066 2638 1246 2677
rect 1066 2604 1067 2638
rect 1101 2604 1139 2638
rect 1173 2604 1211 2638
rect 1245 2604 1246 2638
rect 1066 2565 1246 2604
rect 1066 2531 1067 2565
rect 1101 2531 1139 2565
rect 1173 2531 1211 2565
rect 1245 2531 1246 2565
rect 1066 2492 1246 2531
rect 1066 2458 1067 2492
rect 1101 2482 1139 2492
rect 1101 2458 1103 2482
rect 1066 2448 1103 2458
rect 1137 2458 1139 2482
rect 1173 2482 1211 2492
rect 1173 2458 1175 2482
rect 1137 2448 1175 2458
rect 1209 2458 1211 2482
rect 1245 2458 1246 2492
rect 1209 2448 1246 2458
rect 1066 2419 1246 2448
rect 1066 2385 1067 2419
rect 1101 2414 1139 2419
rect 1101 2385 1103 2414
rect 1066 2380 1103 2385
rect 1137 2385 1139 2414
rect 1173 2414 1211 2419
rect 1173 2385 1175 2414
rect 1137 2380 1175 2385
rect 1209 2385 1211 2414
rect 1245 2385 1246 2419
rect 1209 2380 1246 2385
rect 1066 2346 1246 2380
rect 1066 2312 1067 2346
rect 1101 2312 1103 2346
rect 1137 2312 1139 2346
rect 1173 2312 1175 2346
rect 1209 2312 1211 2346
rect 1245 2312 1246 2346
rect 1066 2278 1246 2312
rect 1066 2273 1103 2278
rect 1066 2239 1067 2273
rect 1101 2244 1103 2273
rect 1137 2273 1175 2278
rect 1137 2244 1139 2273
rect 1101 2239 1139 2244
rect 1173 2244 1175 2273
rect 1209 2273 1246 2278
rect 1209 2244 1211 2273
rect 1173 2239 1211 2244
rect 1245 2239 1246 2273
rect 1066 2210 1246 2239
rect 1066 2200 1103 2210
rect 1066 2166 1067 2200
rect 1101 2176 1103 2200
rect 1137 2200 1175 2210
rect 1137 2176 1139 2200
rect 1101 2166 1139 2176
rect 1173 2176 1175 2200
rect 1209 2200 1246 2210
rect 1209 2176 1211 2200
rect 1173 2166 1211 2176
rect 1245 2166 1246 2200
rect 1066 2142 1246 2166
rect 1066 2126 1103 2142
rect 1066 2092 1067 2126
rect 1101 2108 1103 2126
rect 1137 2126 1175 2142
rect 1137 2108 1139 2126
rect 1101 2092 1139 2108
rect 1173 2108 1175 2126
rect 1209 2126 1246 2142
rect 1209 2108 1211 2126
rect 1173 2092 1211 2108
rect 1245 2092 1246 2126
rect 1066 2074 1246 2092
rect 1066 2052 1103 2074
rect 1066 2018 1067 2052
rect 1101 2040 1103 2052
rect 1137 2052 1175 2074
rect 1137 2040 1139 2052
rect 1101 2018 1139 2040
rect 1173 2040 1175 2052
rect 1209 2052 1246 2074
rect 1209 2040 1211 2052
rect 1173 2018 1211 2040
rect 1245 2018 1246 2052
rect 1066 2006 1246 2018
rect 1066 1978 1103 2006
rect 1066 1944 1067 1978
rect 1101 1972 1103 1978
rect 1137 1978 1175 2006
rect 1137 1972 1139 1978
rect 1101 1944 1139 1972
rect 1173 1972 1175 1978
rect 1209 1978 1246 2006
rect 1209 1972 1211 1978
rect 1173 1944 1211 1972
rect 1245 1944 1246 1978
rect 1066 1938 1246 1944
rect 1066 1904 1103 1938
rect 1137 1904 1175 1938
rect 1209 1904 1246 1938
rect 1066 1870 1067 1904
rect 1101 1870 1139 1904
rect 1173 1870 1211 1904
rect 1245 1870 1246 1904
rect 1066 1836 1103 1870
rect 1137 1836 1175 1870
rect 1209 1836 1246 1870
rect 1066 1830 1246 1836
rect 1066 1796 1067 1830
rect 1101 1802 1139 1830
rect 1101 1796 1103 1802
rect 1066 1768 1103 1796
rect 1137 1796 1139 1802
rect 1173 1802 1211 1830
rect 1173 1796 1175 1802
rect 1137 1768 1175 1796
rect 1209 1796 1211 1802
rect 1245 1796 1246 1830
rect 1209 1768 1246 1796
rect 1066 1756 1246 1768
rect 1066 1722 1067 1756
rect 1101 1734 1139 1756
rect 1101 1722 1103 1734
rect 1066 1700 1103 1722
rect 1137 1722 1139 1734
rect 1173 1734 1211 1756
rect 1173 1722 1175 1734
rect 1137 1700 1175 1722
rect 1209 1722 1211 1734
rect 1245 1722 1246 1756
rect 1209 1700 1246 1722
rect 1066 1682 1246 1700
rect 1066 1648 1067 1682
rect 1101 1666 1139 1682
rect 1101 1648 1103 1666
rect 1066 1632 1103 1648
rect 1137 1648 1139 1666
rect 1173 1666 1211 1682
rect 1173 1648 1175 1666
rect 1137 1632 1175 1648
rect 1209 1648 1211 1666
rect 1245 1648 1246 1682
rect 1209 1632 1246 1648
rect 1066 1608 1246 1632
rect 1066 1574 1067 1608
rect 1101 1598 1139 1608
rect 1101 1574 1103 1598
rect 1066 1564 1103 1574
rect 1137 1574 1139 1598
rect 1173 1598 1211 1608
rect 1173 1574 1175 1598
rect 1137 1564 1175 1574
rect 1209 1574 1211 1598
rect 1245 1574 1246 1608
rect 1209 1564 1246 1574
rect 1066 1548 1246 1564
rect 1311 3104 1431 4200
rect 1873 4308 1993 4324
rect 1873 4274 1916 4308
rect 1950 4274 1993 4308
rect 1873 4234 1993 4274
rect 1873 4200 1916 4234
rect 1950 4200 1993 4234
rect 1311 3070 1354 3104
rect 1388 3070 1431 3104
rect 1311 3026 1431 3070
rect 1311 2992 1354 3026
rect 1388 2992 1431 3026
rect 1311 2948 1431 2992
rect 1311 2914 1354 2948
rect 1388 2914 1431 2948
rect 1311 2870 1431 2914
rect 1311 2836 1354 2870
rect 1388 2836 1431 2870
rect 1311 2792 1431 2836
rect 1311 2758 1354 2792
rect 1388 2758 1431 2792
rect 1311 2713 1431 2758
rect 1311 2679 1354 2713
rect 1388 2679 1431 2713
rect 1311 2634 1431 2679
rect 1311 2600 1354 2634
rect 1388 2600 1431 2634
rect 881 1470 924 1504
rect 958 1470 1001 1504
rect 881 1430 1001 1470
rect 881 1396 924 1430
rect 958 1396 1001 1430
rect 881 1250 1001 1396
rect 881 1216 924 1250
rect 958 1216 1001 1250
rect 881 1178 1001 1216
rect 881 1144 924 1178
rect 958 1144 1001 1178
rect 1311 1504 1431 2600
rect 1533 4092 1635 4118
rect 1669 4092 1771 4118
rect 1533 4082 1563 4092
rect 1741 4082 1771 4092
rect 1533 4014 1563 4048
rect 1741 4014 1771 4048
rect 1533 3946 1563 3980
rect 1741 3946 1771 3980
rect 1533 3878 1563 3912
rect 1741 3878 1771 3912
rect 1533 3810 1563 3844
rect 1741 3810 1771 3844
rect 1533 3742 1563 3776
rect 1741 3742 1771 3776
rect 1533 3674 1563 3708
rect 1741 3674 1771 3708
rect 1533 3606 1563 3640
rect 1741 3606 1771 3640
rect 1533 3538 1563 3572
rect 1741 3538 1771 3572
rect 1533 3470 1563 3504
rect 1741 3470 1771 3504
rect 1533 3402 1563 3436
rect 1741 3402 1771 3436
rect 1533 3334 1563 3368
rect 1741 3334 1771 3368
rect 1533 3266 1563 3300
rect 1741 3266 1771 3300
rect 1533 3198 1563 3232
rect 1741 3198 1771 3232
rect 1567 3164 1635 3194
rect 1669 3164 1737 3194
rect 1533 3148 1635 3164
rect 1669 3148 1771 3164
rect 1533 3108 1771 3148
rect 1533 3074 1563 3108
rect 1597 3074 1635 3108
rect 1669 3074 1707 3108
rect 1741 3074 1771 3108
rect 1533 3044 1771 3074
rect 1533 3028 1601 3044
rect 1533 2994 1563 3028
rect 1597 3010 1601 3028
rect 1635 3028 1669 3044
rect 1597 2994 1635 3010
rect 1703 3028 1771 3044
rect 1703 3010 1707 3028
rect 1669 2994 1707 3010
rect 1741 2994 1771 3028
rect 1533 2974 1771 2994
rect 1533 2948 1601 2974
rect 1533 2914 1563 2948
rect 1597 2940 1601 2948
rect 1635 2948 1669 2974
rect 1597 2914 1635 2940
rect 1703 2948 1771 2974
rect 1703 2940 1707 2948
rect 1669 2914 1707 2940
rect 1741 2914 1771 2948
rect 1533 2904 1771 2914
rect 1533 2870 1601 2904
rect 1635 2870 1669 2904
rect 1703 2870 1771 2904
rect 1533 2868 1771 2870
rect 1533 2834 1563 2868
rect 1597 2834 1635 2868
rect 1669 2834 1707 2868
rect 1741 2834 1771 2868
rect 1533 2800 1601 2834
rect 1635 2800 1669 2834
rect 1703 2800 1771 2834
rect 1533 2788 1771 2800
rect 1533 2754 1563 2788
rect 1597 2764 1635 2788
rect 1597 2754 1601 2764
rect 1533 2730 1601 2754
rect 1669 2764 1707 2788
rect 1635 2730 1669 2754
rect 1703 2754 1707 2764
rect 1741 2754 1771 2788
rect 1703 2730 1771 2754
rect 1533 2708 1771 2730
rect 1533 2674 1563 2708
rect 1597 2694 1635 2708
rect 1597 2674 1601 2694
rect 1533 2660 1601 2674
rect 1669 2694 1707 2708
rect 1635 2660 1669 2674
rect 1703 2674 1707 2694
rect 1741 2674 1771 2708
rect 1703 2660 1771 2674
rect 1533 2628 1771 2660
rect 1533 2594 1563 2628
rect 1597 2594 1635 2628
rect 1669 2594 1707 2628
rect 1741 2594 1771 2628
rect 1533 2556 1771 2594
rect 1533 2540 1635 2556
rect 1669 2540 1771 2556
rect 1567 2518 1635 2540
rect 1669 2518 1737 2540
rect 1533 2472 1563 2506
rect 1741 2472 1771 2506
rect 1533 2404 1563 2438
rect 1741 2404 1771 2438
rect 1533 2336 1563 2370
rect 1741 2336 1771 2370
rect 1533 2268 1563 2302
rect 1741 2268 1771 2302
rect 1533 2200 1563 2234
rect 1741 2200 1771 2234
rect 1533 2132 1563 2166
rect 1741 2132 1771 2166
rect 1533 2064 1563 2098
rect 1741 2064 1771 2098
rect 1533 1996 1563 2030
rect 1741 1996 1771 2030
rect 1533 1928 1563 1962
rect 1741 1928 1771 1962
rect 1533 1860 1563 1894
rect 1741 1860 1771 1894
rect 1533 1792 1563 1826
rect 1741 1792 1771 1826
rect 1533 1724 1563 1758
rect 1741 1724 1771 1758
rect 1533 1656 1563 1690
rect 1741 1656 1771 1690
rect 1533 1620 1563 1622
rect 1741 1620 1771 1622
rect 1533 1586 1635 1620
rect 1669 1586 1771 1620
rect 1533 1536 1771 1586
rect 1873 3104 1993 4200
rect 2303 4308 2423 4324
rect 2303 4274 2346 4308
rect 2380 4274 2423 4308
rect 2303 4234 2423 4274
rect 2303 4200 2346 4234
rect 2380 4200 2423 4234
rect 1873 3070 1916 3104
rect 1950 3070 1993 3104
rect 1873 3026 1993 3070
rect 1873 2992 1916 3026
rect 1950 2992 1993 3026
rect 1873 2948 1993 2992
rect 1873 2914 1916 2948
rect 1950 2914 1993 2948
rect 1873 2870 1993 2914
rect 1873 2836 1916 2870
rect 1950 2836 1993 2870
rect 1873 2792 1993 2836
rect 1873 2758 1916 2792
rect 1950 2758 1993 2792
rect 1873 2713 1993 2758
rect 1873 2679 1916 2713
rect 1950 2679 1993 2713
rect 1873 2634 1993 2679
rect 1873 2600 1916 2634
rect 1950 2600 1993 2634
rect 1311 1470 1354 1504
rect 1388 1470 1431 1504
rect 1311 1430 1431 1470
rect 1311 1396 1354 1430
rect 1388 1396 1431 1430
rect 1311 1250 1431 1396
rect 1311 1144 1318 1250
rect 1424 1144 1431 1250
rect 1873 1504 1993 2600
rect 2058 4064 2059 4098
rect 2093 4082 2131 4098
rect 2093 4064 2095 4082
rect 2058 4048 2095 4064
rect 2129 4064 2131 4082
rect 2165 4082 2203 4098
rect 2165 4064 2167 4082
rect 2129 4048 2167 4064
rect 2201 4064 2203 4082
rect 2237 4064 2238 4098
rect 2201 4048 2238 4064
rect 2058 4025 2238 4048
rect 2058 3991 2059 4025
rect 2093 4014 2131 4025
rect 2093 3991 2095 4014
rect 2058 3980 2095 3991
rect 2129 3991 2131 4014
rect 2165 4014 2203 4025
rect 2165 3991 2167 4014
rect 2129 3980 2167 3991
rect 2201 3991 2203 4014
rect 2237 3991 2238 4025
rect 2201 3980 2238 3991
rect 2058 3952 2238 3980
rect 2058 3918 2059 3952
rect 2093 3946 2131 3952
rect 2093 3918 2095 3946
rect 2058 3912 2095 3918
rect 2129 3918 2131 3946
rect 2165 3946 2203 3952
rect 2165 3918 2167 3946
rect 2129 3912 2167 3918
rect 2201 3918 2203 3946
rect 2237 3918 2238 3952
rect 2201 3912 2238 3918
rect 2058 3879 2238 3912
rect 2058 3845 2059 3879
rect 2093 3878 2131 3879
rect 2093 3845 2095 3878
rect 2058 3844 2095 3845
rect 2129 3845 2131 3878
rect 2165 3878 2203 3879
rect 2165 3845 2167 3878
rect 2129 3844 2167 3845
rect 2201 3845 2203 3878
rect 2237 3845 2238 3879
rect 2201 3844 2238 3845
rect 2058 3810 2238 3844
rect 2058 3806 2095 3810
rect 2058 3772 2059 3806
rect 2093 3776 2095 3806
rect 2129 3806 2167 3810
rect 2129 3776 2131 3806
rect 2093 3772 2131 3776
rect 2165 3776 2167 3806
rect 2201 3806 2238 3810
rect 2201 3776 2203 3806
rect 2165 3772 2203 3776
rect 2237 3772 2238 3806
rect 2058 3742 2238 3772
rect 2058 3733 2095 3742
rect 2058 3699 2059 3733
rect 2093 3708 2095 3733
rect 2129 3733 2167 3742
rect 2129 3708 2131 3733
rect 2093 3699 2131 3708
rect 2165 3708 2167 3733
rect 2201 3733 2238 3742
rect 2201 3708 2203 3733
rect 2165 3699 2203 3708
rect 2237 3699 2238 3733
rect 2058 3674 2238 3699
rect 2058 3660 2095 3674
rect 2058 3626 2059 3660
rect 2093 3640 2095 3660
rect 2129 3660 2167 3674
rect 2129 3640 2131 3660
rect 2093 3626 2131 3640
rect 2165 3640 2167 3660
rect 2201 3660 2238 3674
rect 2201 3640 2203 3660
rect 2165 3626 2203 3640
rect 2237 3626 2238 3660
rect 2058 3606 2238 3626
rect 2058 3587 2095 3606
rect 2058 3553 2059 3587
rect 2093 3572 2095 3587
rect 2129 3587 2167 3606
rect 2129 3572 2131 3587
rect 2093 3553 2131 3572
rect 2165 3572 2167 3587
rect 2201 3587 2238 3606
rect 2201 3572 2203 3587
rect 2165 3553 2203 3572
rect 2237 3553 2238 3587
rect 2058 3538 2238 3553
rect 2058 3514 2095 3538
rect 2058 3480 2059 3514
rect 2093 3504 2095 3514
rect 2129 3514 2167 3538
rect 2129 3504 2131 3514
rect 2093 3480 2131 3504
rect 2165 3504 2167 3514
rect 2201 3514 2238 3538
rect 2201 3504 2203 3514
rect 2165 3480 2203 3504
rect 2237 3480 2238 3514
rect 2058 3470 2238 3480
rect 2058 3441 2095 3470
rect 2058 3407 2059 3441
rect 2093 3436 2095 3441
rect 2129 3441 2167 3470
rect 2129 3436 2131 3441
rect 2093 3407 2131 3436
rect 2165 3436 2167 3441
rect 2201 3441 2238 3470
rect 2201 3436 2203 3441
rect 2165 3407 2203 3436
rect 2237 3407 2238 3441
rect 2058 3402 2238 3407
rect 2058 3368 2095 3402
rect 2129 3368 2167 3402
rect 2201 3368 2238 3402
rect 2058 3334 2059 3368
rect 2093 3334 2131 3368
rect 2165 3334 2203 3368
rect 2237 3334 2238 3368
rect 2058 3300 2095 3334
rect 2129 3300 2167 3334
rect 2201 3300 2238 3334
rect 2058 3295 2238 3300
rect 2058 3261 2059 3295
rect 2093 3266 2131 3295
rect 2093 3261 2095 3266
rect 2058 3232 2095 3261
rect 2129 3261 2131 3266
rect 2165 3266 2203 3295
rect 2165 3261 2167 3266
rect 2129 3232 2167 3261
rect 2201 3261 2203 3266
rect 2237 3261 2238 3295
rect 2201 3232 2238 3261
rect 2058 3222 2238 3232
rect 2058 3188 2059 3222
rect 2093 3198 2131 3222
rect 2093 3188 2095 3198
rect 2058 3164 2095 3188
rect 2129 3188 2131 3198
rect 2165 3198 2203 3222
rect 2165 3188 2167 3198
rect 2129 3164 2167 3188
rect 2201 3188 2203 3198
rect 2237 3188 2238 3222
rect 2201 3164 2238 3188
rect 2058 3149 2238 3164
rect 2058 3115 2059 3149
rect 2093 3115 2131 3149
rect 2165 3115 2203 3149
rect 2237 3115 2238 3149
rect 2058 3076 2238 3115
rect 2058 3042 2059 3076
rect 2093 3042 2131 3076
rect 2165 3042 2203 3076
rect 2237 3042 2238 3076
rect 2058 3003 2238 3042
rect 2058 2969 2059 3003
rect 2093 2969 2131 3003
rect 2165 2969 2203 3003
rect 2237 2969 2238 3003
rect 2058 2930 2238 2969
rect 2058 2896 2059 2930
rect 2093 2896 2131 2930
rect 2165 2896 2203 2930
rect 2237 2896 2238 2930
rect 2058 2857 2238 2896
rect 2058 2823 2059 2857
rect 2093 2823 2131 2857
rect 2165 2823 2203 2857
rect 2237 2823 2238 2857
rect 2058 2784 2238 2823
rect 2058 2750 2059 2784
rect 2093 2750 2131 2784
rect 2165 2750 2203 2784
rect 2237 2750 2238 2784
rect 2058 2711 2238 2750
rect 2058 2677 2059 2711
rect 2093 2677 2131 2711
rect 2165 2677 2203 2711
rect 2237 2677 2238 2711
rect 2058 2638 2238 2677
rect 2058 2604 2059 2638
rect 2093 2604 2131 2638
rect 2165 2604 2203 2638
rect 2237 2604 2238 2638
rect 2058 2565 2238 2604
rect 2058 2531 2059 2565
rect 2093 2531 2131 2565
rect 2165 2531 2203 2565
rect 2237 2531 2238 2565
rect 2058 2492 2238 2531
rect 2058 2458 2059 2492
rect 2093 2482 2131 2492
rect 2093 2458 2095 2482
rect 2058 2448 2095 2458
rect 2129 2458 2131 2482
rect 2165 2482 2203 2492
rect 2165 2458 2167 2482
rect 2129 2448 2167 2458
rect 2201 2458 2203 2482
rect 2237 2458 2238 2492
rect 2201 2448 2238 2458
rect 2058 2419 2238 2448
rect 2058 2385 2059 2419
rect 2093 2414 2131 2419
rect 2093 2385 2095 2414
rect 2058 2380 2095 2385
rect 2129 2385 2131 2414
rect 2165 2414 2203 2419
rect 2165 2385 2167 2414
rect 2129 2380 2167 2385
rect 2201 2385 2203 2414
rect 2237 2385 2238 2419
rect 2201 2380 2238 2385
rect 2058 2346 2238 2380
rect 2058 2312 2059 2346
rect 2093 2312 2095 2346
rect 2129 2312 2131 2346
rect 2165 2312 2167 2346
rect 2201 2312 2203 2346
rect 2237 2312 2238 2346
rect 2058 2278 2238 2312
rect 2058 2273 2095 2278
rect 2058 2239 2059 2273
rect 2093 2244 2095 2273
rect 2129 2273 2167 2278
rect 2129 2244 2131 2273
rect 2093 2239 2131 2244
rect 2165 2244 2167 2273
rect 2201 2273 2238 2278
rect 2201 2244 2203 2273
rect 2165 2239 2203 2244
rect 2237 2239 2238 2273
rect 2058 2210 2238 2239
rect 2058 2200 2095 2210
rect 2058 2166 2059 2200
rect 2093 2176 2095 2200
rect 2129 2200 2167 2210
rect 2129 2176 2131 2200
rect 2093 2166 2131 2176
rect 2165 2176 2167 2200
rect 2201 2200 2238 2210
rect 2201 2176 2203 2200
rect 2165 2166 2203 2176
rect 2237 2166 2238 2200
rect 2058 2142 2238 2166
rect 2058 2126 2095 2142
rect 2058 2092 2059 2126
rect 2093 2108 2095 2126
rect 2129 2126 2167 2142
rect 2129 2108 2131 2126
rect 2093 2092 2131 2108
rect 2165 2108 2167 2126
rect 2201 2126 2238 2142
rect 2201 2108 2203 2126
rect 2165 2092 2203 2108
rect 2237 2092 2238 2126
rect 2058 2074 2238 2092
rect 2058 2052 2095 2074
rect 2058 2018 2059 2052
rect 2093 2040 2095 2052
rect 2129 2052 2167 2074
rect 2129 2040 2131 2052
rect 2093 2018 2131 2040
rect 2165 2040 2167 2052
rect 2201 2052 2238 2074
rect 2201 2040 2203 2052
rect 2165 2018 2203 2040
rect 2237 2018 2238 2052
rect 2058 2006 2238 2018
rect 2058 1978 2095 2006
rect 2058 1944 2059 1978
rect 2093 1972 2095 1978
rect 2129 1978 2167 2006
rect 2129 1972 2131 1978
rect 2093 1944 2131 1972
rect 2165 1972 2167 1978
rect 2201 1978 2238 2006
rect 2201 1972 2203 1978
rect 2165 1944 2203 1972
rect 2237 1944 2238 1978
rect 2058 1938 2238 1944
rect 2058 1904 2095 1938
rect 2129 1904 2167 1938
rect 2201 1904 2238 1938
rect 2058 1870 2059 1904
rect 2093 1870 2131 1904
rect 2165 1870 2203 1904
rect 2237 1870 2238 1904
rect 2058 1836 2095 1870
rect 2129 1836 2167 1870
rect 2201 1836 2238 1870
rect 2058 1830 2238 1836
rect 2058 1796 2059 1830
rect 2093 1802 2131 1830
rect 2093 1796 2095 1802
rect 2058 1768 2095 1796
rect 2129 1796 2131 1802
rect 2165 1802 2203 1830
rect 2165 1796 2167 1802
rect 2129 1768 2167 1796
rect 2201 1796 2203 1802
rect 2237 1796 2238 1830
rect 2201 1768 2238 1796
rect 2058 1756 2238 1768
rect 2058 1722 2059 1756
rect 2093 1734 2131 1756
rect 2093 1722 2095 1734
rect 2058 1700 2095 1722
rect 2129 1722 2131 1734
rect 2165 1734 2203 1756
rect 2165 1722 2167 1734
rect 2129 1700 2167 1722
rect 2201 1722 2203 1734
rect 2237 1722 2238 1756
rect 2201 1700 2238 1722
rect 2058 1682 2238 1700
rect 2058 1648 2059 1682
rect 2093 1666 2131 1682
rect 2093 1648 2095 1666
rect 2058 1632 2095 1648
rect 2129 1648 2131 1666
rect 2165 1666 2203 1682
rect 2165 1648 2167 1666
rect 2129 1632 2167 1648
rect 2201 1648 2203 1666
rect 2237 1648 2238 1682
rect 2201 1632 2238 1648
rect 2058 1608 2238 1632
rect 2058 1574 2059 1608
rect 2093 1598 2131 1608
rect 2093 1574 2095 1598
rect 2058 1564 2095 1574
rect 2129 1574 2131 1598
rect 2165 1598 2203 1608
rect 2165 1574 2167 1598
rect 2129 1564 2167 1574
rect 2201 1574 2203 1598
rect 2237 1574 2238 1608
rect 2201 1564 2238 1574
rect 2058 1548 2238 1564
rect 2303 3104 2423 4200
rect 2865 4308 2985 4324
rect 2865 4274 2908 4308
rect 2942 4274 2985 4308
rect 2865 4234 2985 4274
rect 2865 4200 2908 4234
rect 2942 4200 2985 4234
rect 2303 3070 2346 3104
rect 2380 3070 2423 3104
rect 2303 3026 2423 3070
rect 2303 2992 2346 3026
rect 2380 2992 2423 3026
rect 2303 2948 2423 2992
rect 2303 2914 2346 2948
rect 2380 2914 2423 2948
rect 2303 2870 2423 2914
rect 2303 2836 2346 2870
rect 2380 2836 2423 2870
rect 2303 2792 2423 2836
rect 2303 2758 2346 2792
rect 2380 2758 2423 2792
rect 2303 2713 2423 2758
rect 2303 2679 2346 2713
rect 2380 2679 2423 2713
rect 2303 2634 2423 2679
rect 2303 2600 2346 2634
rect 2380 2600 2423 2634
rect 1873 1470 1916 1504
rect 1950 1470 1993 1504
rect 1873 1430 1993 1470
rect 1873 1396 1916 1430
rect 1950 1396 1993 1430
rect 1873 1250 1993 1396
rect 1873 1144 1880 1250
rect 1986 1144 1993 1250
rect 2303 1504 2423 2600
rect 2525 4092 2627 4118
rect 2661 4092 2763 4118
rect 2525 4082 2555 4092
rect 2733 4082 2763 4092
rect 2525 4014 2555 4048
rect 2733 4014 2763 4048
rect 2525 3946 2555 3980
rect 2733 3946 2763 3980
rect 2525 3878 2555 3912
rect 2733 3878 2763 3912
rect 2525 3810 2555 3844
rect 2733 3810 2763 3844
rect 2525 3742 2555 3776
rect 2733 3742 2763 3776
rect 2525 3674 2555 3708
rect 2733 3674 2763 3708
rect 2525 3606 2555 3640
rect 2733 3606 2763 3640
rect 2525 3538 2555 3572
rect 2733 3538 2763 3572
rect 2525 3470 2555 3504
rect 2733 3470 2763 3504
rect 2525 3402 2555 3436
rect 2733 3402 2763 3436
rect 2525 3334 2555 3368
rect 2733 3334 2763 3368
rect 2525 3266 2555 3300
rect 2733 3266 2763 3300
rect 2525 3198 2555 3232
rect 2733 3198 2763 3232
rect 2559 3164 2627 3194
rect 2661 3164 2729 3194
rect 2525 3148 2627 3164
rect 2661 3148 2763 3164
rect 2525 3108 2763 3148
rect 2525 3074 2555 3108
rect 2589 3074 2627 3108
rect 2661 3074 2699 3108
rect 2733 3074 2763 3108
rect 2525 3044 2763 3074
rect 2525 3028 2593 3044
rect 2525 2994 2555 3028
rect 2589 3010 2593 3028
rect 2627 3028 2661 3044
rect 2589 2994 2627 3010
rect 2695 3028 2763 3044
rect 2695 3010 2699 3028
rect 2661 2994 2699 3010
rect 2733 2994 2763 3028
rect 2525 2974 2763 2994
rect 2525 2948 2593 2974
rect 2525 2914 2555 2948
rect 2589 2940 2593 2948
rect 2627 2948 2661 2974
rect 2589 2914 2627 2940
rect 2695 2948 2763 2974
rect 2695 2940 2699 2948
rect 2661 2914 2699 2940
rect 2733 2914 2763 2948
rect 2525 2904 2763 2914
rect 2525 2870 2593 2904
rect 2627 2870 2661 2904
rect 2695 2870 2763 2904
rect 2525 2868 2763 2870
rect 2525 2834 2555 2868
rect 2589 2834 2627 2868
rect 2661 2834 2699 2868
rect 2733 2834 2763 2868
rect 2525 2800 2593 2834
rect 2627 2800 2661 2834
rect 2695 2800 2763 2834
rect 2525 2788 2763 2800
rect 2525 2754 2555 2788
rect 2589 2764 2627 2788
rect 2589 2754 2593 2764
rect 2525 2730 2593 2754
rect 2661 2764 2699 2788
rect 2627 2730 2661 2754
rect 2695 2754 2699 2764
rect 2733 2754 2763 2788
rect 2695 2730 2763 2754
rect 2525 2708 2763 2730
rect 2525 2674 2555 2708
rect 2589 2694 2627 2708
rect 2589 2674 2593 2694
rect 2525 2660 2593 2674
rect 2661 2694 2699 2708
rect 2627 2660 2661 2674
rect 2695 2674 2699 2694
rect 2733 2674 2763 2708
rect 2695 2660 2763 2674
rect 2525 2628 2763 2660
rect 2525 2594 2555 2628
rect 2589 2594 2627 2628
rect 2661 2594 2699 2628
rect 2733 2594 2763 2628
rect 2525 2556 2763 2594
rect 2525 2540 2627 2556
rect 2661 2540 2763 2556
rect 2559 2518 2627 2540
rect 2661 2518 2729 2540
rect 2525 2472 2555 2506
rect 2733 2472 2763 2506
rect 2525 2404 2555 2438
rect 2733 2404 2763 2438
rect 2525 2336 2555 2370
rect 2733 2336 2763 2370
rect 2525 2268 2555 2302
rect 2733 2268 2763 2302
rect 2525 2200 2555 2234
rect 2733 2200 2763 2234
rect 2525 2132 2555 2166
rect 2733 2132 2763 2166
rect 2525 2064 2555 2098
rect 2733 2064 2763 2098
rect 2525 1996 2555 2030
rect 2733 1996 2763 2030
rect 2525 1928 2555 1962
rect 2733 1928 2763 1962
rect 2525 1860 2555 1894
rect 2733 1860 2763 1894
rect 2525 1792 2555 1826
rect 2733 1792 2763 1826
rect 2525 1724 2555 1758
rect 2733 1724 2763 1758
rect 2525 1656 2555 1690
rect 2733 1656 2763 1690
rect 2525 1620 2555 1622
rect 2733 1620 2763 1622
rect 2525 1586 2627 1620
rect 2661 1586 2763 1620
rect 2525 1536 2763 1586
rect 2865 3104 2985 4200
rect 3295 4308 3415 4324
rect 3295 4274 3338 4308
rect 3372 4274 3415 4308
rect 3295 4234 3415 4274
rect 3295 4200 3338 4234
rect 3372 4200 3415 4234
rect 2865 3070 2908 3104
rect 2942 3070 2985 3104
rect 2865 3026 2985 3070
rect 2865 2992 2908 3026
rect 2942 2992 2985 3026
rect 2865 2948 2985 2992
rect 2865 2914 2908 2948
rect 2942 2914 2985 2948
rect 2865 2870 2985 2914
rect 2865 2836 2908 2870
rect 2942 2836 2985 2870
rect 2865 2792 2985 2836
rect 2865 2758 2908 2792
rect 2942 2758 2985 2792
rect 2865 2713 2985 2758
rect 2865 2679 2908 2713
rect 2942 2679 2985 2713
rect 2865 2634 2985 2679
rect 2865 2600 2908 2634
rect 2942 2600 2985 2634
rect 2303 1470 2346 1504
rect 2380 1470 2423 1504
rect 2303 1430 2423 1470
rect 2303 1396 2346 1430
rect 2380 1396 2423 1430
rect 2303 1250 2423 1396
rect 2303 1144 2310 1250
rect 2416 1144 2423 1250
rect 2865 1504 2985 2600
rect 3050 4064 3051 4098
rect 3085 4082 3123 4098
rect 3085 4064 3087 4082
rect 3050 4048 3087 4064
rect 3121 4064 3123 4082
rect 3157 4082 3195 4098
rect 3157 4064 3159 4082
rect 3121 4048 3159 4064
rect 3193 4064 3195 4082
rect 3229 4064 3230 4098
rect 3193 4048 3230 4064
rect 3050 4025 3230 4048
rect 3050 3991 3051 4025
rect 3085 4014 3123 4025
rect 3085 3991 3087 4014
rect 3050 3980 3087 3991
rect 3121 3991 3123 4014
rect 3157 4014 3195 4025
rect 3157 3991 3159 4014
rect 3121 3980 3159 3991
rect 3193 3991 3195 4014
rect 3229 3991 3230 4025
rect 3193 3980 3230 3991
rect 3050 3952 3230 3980
rect 3050 3918 3051 3952
rect 3085 3946 3123 3952
rect 3085 3918 3087 3946
rect 3050 3912 3087 3918
rect 3121 3918 3123 3946
rect 3157 3946 3195 3952
rect 3157 3918 3159 3946
rect 3121 3912 3159 3918
rect 3193 3918 3195 3946
rect 3229 3918 3230 3952
rect 3193 3912 3230 3918
rect 3050 3879 3230 3912
rect 3050 3845 3051 3879
rect 3085 3878 3123 3879
rect 3085 3845 3087 3878
rect 3050 3844 3087 3845
rect 3121 3845 3123 3878
rect 3157 3878 3195 3879
rect 3157 3845 3159 3878
rect 3121 3844 3159 3845
rect 3193 3845 3195 3878
rect 3229 3845 3230 3879
rect 3193 3844 3230 3845
rect 3050 3810 3230 3844
rect 3050 3806 3087 3810
rect 3050 3772 3051 3806
rect 3085 3776 3087 3806
rect 3121 3806 3159 3810
rect 3121 3776 3123 3806
rect 3085 3772 3123 3776
rect 3157 3776 3159 3806
rect 3193 3806 3230 3810
rect 3193 3776 3195 3806
rect 3157 3772 3195 3776
rect 3229 3772 3230 3806
rect 3050 3742 3230 3772
rect 3050 3733 3087 3742
rect 3050 3699 3051 3733
rect 3085 3708 3087 3733
rect 3121 3733 3159 3742
rect 3121 3708 3123 3733
rect 3085 3699 3123 3708
rect 3157 3708 3159 3733
rect 3193 3733 3230 3742
rect 3193 3708 3195 3733
rect 3157 3699 3195 3708
rect 3229 3699 3230 3733
rect 3050 3674 3230 3699
rect 3050 3660 3087 3674
rect 3050 3626 3051 3660
rect 3085 3640 3087 3660
rect 3121 3660 3159 3674
rect 3121 3640 3123 3660
rect 3085 3626 3123 3640
rect 3157 3640 3159 3660
rect 3193 3660 3230 3674
rect 3193 3640 3195 3660
rect 3157 3626 3195 3640
rect 3229 3626 3230 3660
rect 3050 3606 3230 3626
rect 3050 3587 3087 3606
rect 3050 3553 3051 3587
rect 3085 3572 3087 3587
rect 3121 3587 3159 3606
rect 3121 3572 3123 3587
rect 3085 3553 3123 3572
rect 3157 3572 3159 3587
rect 3193 3587 3230 3606
rect 3193 3572 3195 3587
rect 3157 3553 3195 3572
rect 3229 3553 3230 3587
rect 3050 3538 3230 3553
rect 3050 3514 3087 3538
rect 3050 3480 3051 3514
rect 3085 3504 3087 3514
rect 3121 3514 3159 3538
rect 3121 3504 3123 3514
rect 3085 3480 3123 3504
rect 3157 3504 3159 3514
rect 3193 3514 3230 3538
rect 3193 3504 3195 3514
rect 3157 3480 3195 3504
rect 3229 3480 3230 3514
rect 3050 3470 3230 3480
rect 3050 3441 3087 3470
rect 3050 3407 3051 3441
rect 3085 3436 3087 3441
rect 3121 3441 3159 3470
rect 3121 3436 3123 3441
rect 3085 3407 3123 3436
rect 3157 3436 3159 3441
rect 3193 3441 3230 3470
rect 3193 3436 3195 3441
rect 3157 3407 3195 3436
rect 3229 3407 3230 3441
rect 3050 3402 3230 3407
rect 3050 3368 3087 3402
rect 3121 3368 3159 3402
rect 3193 3368 3230 3402
rect 3050 3334 3051 3368
rect 3085 3334 3123 3368
rect 3157 3334 3195 3368
rect 3229 3334 3230 3368
rect 3050 3300 3087 3334
rect 3121 3300 3159 3334
rect 3193 3300 3230 3334
rect 3050 3295 3230 3300
rect 3050 3261 3051 3295
rect 3085 3266 3123 3295
rect 3085 3261 3087 3266
rect 3050 3232 3087 3261
rect 3121 3261 3123 3266
rect 3157 3266 3195 3295
rect 3157 3261 3159 3266
rect 3121 3232 3159 3261
rect 3193 3261 3195 3266
rect 3229 3261 3230 3295
rect 3193 3232 3230 3261
rect 3050 3222 3230 3232
rect 3050 3188 3051 3222
rect 3085 3198 3123 3222
rect 3085 3188 3087 3198
rect 3050 3164 3087 3188
rect 3121 3188 3123 3198
rect 3157 3198 3195 3222
rect 3157 3188 3159 3198
rect 3121 3164 3159 3188
rect 3193 3188 3195 3198
rect 3229 3188 3230 3222
rect 3193 3164 3230 3188
rect 3050 3149 3230 3164
rect 3050 3115 3051 3149
rect 3085 3115 3123 3149
rect 3157 3115 3195 3149
rect 3229 3115 3230 3149
rect 3050 3076 3230 3115
rect 3050 3042 3051 3076
rect 3085 3042 3123 3076
rect 3157 3042 3195 3076
rect 3229 3042 3230 3076
rect 3050 3003 3230 3042
rect 3050 2969 3051 3003
rect 3085 2969 3123 3003
rect 3157 2969 3195 3003
rect 3229 2969 3230 3003
rect 3050 2930 3230 2969
rect 3050 2896 3051 2930
rect 3085 2896 3123 2930
rect 3157 2896 3195 2930
rect 3229 2896 3230 2930
rect 3050 2857 3230 2896
rect 3050 2823 3051 2857
rect 3085 2823 3123 2857
rect 3157 2823 3195 2857
rect 3229 2823 3230 2857
rect 3050 2784 3230 2823
rect 3050 2750 3051 2784
rect 3085 2750 3123 2784
rect 3157 2750 3195 2784
rect 3229 2750 3230 2784
rect 3050 2711 3230 2750
rect 3050 2677 3051 2711
rect 3085 2677 3123 2711
rect 3157 2677 3195 2711
rect 3229 2677 3230 2711
rect 3050 2638 3230 2677
rect 3050 2604 3051 2638
rect 3085 2604 3123 2638
rect 3157 2604 3195 2638
rect 3229 2604 3230 2638
rect 3050 2565 3230 2604
rect 3050 2531 3051 2565
rect 3085 2531 3123 2565
rect 3157 2531 3195 2565
rect 3229 2531 3230 2565
rect 3050 2492 3230 2531
rect 3050 2458 3051 2492
rect 3085 2482 3123 2492
rect 3085 2458 3087 2482
rect 3050 2448 3087 2458
rect 3121 2458 3123 2482
rect 3157 2482 3195 2492
rect 3157 2458 3159 2482
rect 3121 2448 3159 2458
rect 3193 2458 3195 2482
rect 3229 2458 3230 2492
rect 3193 2448 3230 2458
rect 3050 2419 3230 2448
rect 3050 2385 3051 2419
rect 3085 2414 3123 2419
rect 3085 2385 3087 2414
rect 3050 2380 3087 2385
rect 3121 2385 3123 2414
rect 3157 2414 3195 2419
rect 3157 2385 3159 2414
rect 3121 2380 3159 2385
rect 3193 2385 3195 2414
rect 3229 2385 3230 2419
rect 3193 2380 3230 2385
rect 3050 2346 3230 2380
rect 3050 2312 3051 2346
rect 3085 2312 3087 2346
rect 3121 2312 3123 2346
rect 3157 2312 3159 2346
rect 3193 2312 3195 2346
rect 3229 2312 3230 2346
rect 3050 2278 3230 2312
rect 3050 2273 3087 2278
rect 3050 2239 3051 2273
rect 3085 2244 3087 2273
rect 3121 2273 3159 2278
rect 3121 2244 3123 2273
rect 3085 2239 3123 2244
rect 3157 2244 3159 2273
rect 3193 2273 3230 2278
rect 3193 2244 3195 2273
rect 3157 2239 3195 2244
rect 3229 2239 3230 2273
rect 3050 2210 3230 2239
rect 3050 2200 3087 2210
rect 3050 2166 3051 2200
rect 3085 2176 3087 2200
rect 3121 2200 3159 2210
rect 3121 2176 3123 2200
rect 3085 2166 3123 2176
rect 3157 2176 3159 2200
rect 3193 2200 3230 2210
rect 3193 2176 3195 2200
rect 3157 2166 3195 2176
rect 3229 2166 3230 2200
rect 3050 2142 3230 2166
rect 3050 2126 3087 2142
rect 3050 2092 3051 2126
rect 3085 2108 3087 2126
rect 3121 2126 3159 2142
rect 3121 2108 3123 2126
rect 3085 2092 3123 2108
rect 3157 2108 3159 2126
rect 3193 2126 3230 2142
rect 3193 2108 3195 2126
rect 3157 2092 3195 2108
rect 3229 2092 3230 2126
rect 3050 2074 3230 2092
rect 3050 2052 3087 2074
rect 3050 2018 3051 2052
rect 3085 2040 3087 2052
rect 3121 2052 3159 2074
rect 3121 2040 3123 2052
rect 3085 2018 3123 2040
rect 3157 2040 3159 2052
rect 3193 2052 3230 2074
rect 3193 2040 3195 2052
rect 3157 2018 3195 2040
rect 3229 2018 3230 2052
rect 3050 2006 3230 2018
rect 3050 1978 3087 2006
rect 3050 1944 3051 1978
rect 3085 1972 3087 1978
rect 3121 1978 3159 2006
rect 3121 1972 3123 1978
rect 3085 1944 3123 1972
rect 3157 1972 3159 1978
rect 3193 1978 3230 2006
rect 3193 1972 3195 1978
rect 3157 1944 3195 1972
rect 3229 1944 3230 1978
rect 3050 1938 3230 1944
rect 3050 1904 3087 1938
rect 3121 1904 3159 1938
rect 3193 1904 3230 1938
rect 3050 1870 3051 1904
rect 3085 1870 3123 1904
rect 3157 1870 3195 1904
rect 3229 1870 3230 1904
rect 3050 1836 3087 1870
rect 3121 1836 3159 1870
rect 3193 1836 3230 1870
rect 3050 1830 3230 1836
rect 3050 1796 3051 1830
rect 3085 1802 3123 1830
rect 3085 1796 3087 1802
rect 3050 1768 3087 1796
rect 3121 1796 3123 1802
rect 3157 1802 3195 1830
rect 3157 1796 3159 1802
rect 3121 1768 3159 1796
rect 3193 1796 3195 1802
rect 3229 1796 3230 1830
rect 3193 1768 3230 1796
rect 3050 1756 3230 1768
rect 3050 1722 3051 1756
rect 3085 1734 3123 1756
rect 3085 1722 3087 1734
rect 3050 1700 3087 1722
rect 3121 1722 3123 1734
rect 3157 1734 3195 1756
rect 3157 1722 3159 1734
rect 3121 1700 3159 1722
rect 3193 1722 3195 1734
rect 3229 1722 3230 1756
rect 3193 1700 3230 1722
rect 3050 1682 3230 1700
rect 3050 1648 3051 1682
rect 3085 1666 3123 1682
rect 3085 1648 3087 1666
rect 3050 1632 3087 1648
rect 3121 1648 3123 1666
rect 3157 1666 3195 1682
rect 3157 1648 3159 1666
rect 3121 1632 3159 1648
rect 3193 1648 3195 1666
rect 3229 1648 3230 1682
rect 3193 1632 3230 1648
rect 3050 1608 3230 1632
rect 3050 1574 3051 1608
rect 3085 1598 3123 1608
rect 3085 1574 3087 1598
rect 3050 1564 3087 1574
rect 3121 1574 3123 1598
rect 3157 1598 3195 1608
rect 3157 1574 3159 1598
rect 3121 1564 3159 1574
rect 3193 1574 3195 1598
rect 3229 1574 3230 1608
rect 3193 1564 3230 1574
rect 3050 1548 3230 1564
rect 3295 3104 3415 4200
rect 3857 4308 3977 4324
rect 3857 4274 3900 4308
rect 3934 4274 3977 4308
rect 3857 4234 3977 4274
rect 3857 4200 3900 4234
rect 3934 4200 3977 4234
rect 3295 3070 3338 3104
rect 3372 3070 3415 3104
rect 3295 3026 3415 3070
rect 3295 2992 3338 3026
rect 3372 2992 3415 3026
rect 3295 2948 3415 2992
rect 3295 2914 3338 2948
rect 3372 2914 3415 2948
rect 3295 2870 3415 2914
rect 3295 2836 3338 2870
rect 3372 2836 3415 2870
rect 3295 2792 3415 2836
rect 3295 2758 3338 2792
rect 3372 2758 3415 2792
rect 3295 2713 3415 2758
rect 3295 2679 3338 2713
rect 3372 2679 3415 2713
rect 3295 2634 3415 2679
rect 3295 2600 3338 2634
rect 3372 2600 3415 2634
rect 2865 1470 2908 1504
rect 2942 1470 2985 1504
rect 2865 1430 2985 1470
rect 2865 1396 2908 1430
rect 2942 1396 2985 1430
rect 2865 1250 2985 1396
rect 2865 1144 2872 1250
rect 2978 1144 2985 1250
rect 3295 1504 3415 2600
rect 3517 4092 3619 4118
rect 3653 4092 3755 4118
rect 3517 4082 3547 4092
rect 3725 4082 3755 4092
rect 3517 4014 3547 4048
rect 3725 4014 3755 4048
rect 3517 3946 3547 3980
rect 3725 3946 3755 3980
rect 3517 3878 3547 3912
rect 3725 3878 3755 3912
rect 3517 3810 3547 3844
rect 3725 3810 3755 3844
rect 3517 3742 3547 3776
rect 3725 3742 3755 3776
rect 3517 3674 3547 3708
rect 3725 3674 3755 3708
rect 3517 3606 3547 3640
rect 3725 3606 3755 3640
rect 3517 3538 3547 3572
rect 3725 3538 3755 3572
rect 3517 3470 3547 3504
rect 3725 3470 3755 3504
rect 3517 3402 3547 3436
rect 3725 3402 3755 3436
rect 3517 3334 3547 3368
rect 3725 3334 3755 3368
rect 3517 3266 3547 3300
rect 3725 3266 3755 3300
rect 3517 3198 3547 3232
rect 3725 3198 3755 3232
rect 3551 3164 3619 3194
rect 3653 3164 3721 3194
rect 3517 3148 3619 3164
rect 3653 3148 3755 3164
rect 3517 3108 3755 3148
rect 3517 3074 3547 3108
rect 3581 3074 3619 3108
rect 3653 3074 3691 3108
rect 3725 3074 3755 3108
rect 3517 3044 3755 3074
rect 3517 3028 3585 3044
rect 3517 2994 3547 3028
rect 3581 3010 3585 3028
rect 3619 3028 3653 3044
rect 3581 2994 3619 3010
rect 3687 3028 3755 3044
rect 3687 3010 3691 3028
rect 3653 2994 3691 3010
rect 3725 2994 3755 3028
rect 3517 2974 3755 2994
rect 3517 2948 3585 2974
rect 3517 2914 3547 2948
rect 3581 2940 3585 2948
rect 3619 2948 3653 2974
rect 3581 2914 3619 2940
rect 3687 2948 3755 2974
rect 3687 2940 3691 2948
rect 3653 2914 3691 2940
rect 3725 2914 3755 2948
rect 3517 2904 3755 2914
rect 3517 2870 3585 2904
rect 3619 2870 3653 2904
rect 3687 2870 3755 2904
rect 3517 2868 3755 2870
rect 3517 2834 3547 2868
rect 3581 2834 3619 2868
rect 3653 2834 3691 2868
rect 3725 2834 3755 2868
rect 3517 2800 3585 2834
rect 3619 2800 3653 2834
rect 3687 2800 3755 2834
rect 3517 2788 3755 2800
rect 3517 2754 3547 2788
rect 3581 2764 3619 2788
rect 3581 2754 3585 2764
rect 3517 2730 3585 2754
rect 3653 2764 3691 2788
rect 3619 2730 3653 2754
rect 3687 2754 3691 2764
rect 3725 2754 3755 2788
rect 3687 2730 3755 2754
rect 3517 2708 3755 2730
rect 3517 2674 3547 2708
rect 3581 2694 3619 2708
rect 3581 2674 3585 2694
rect 3517 2660 3585 2674
rect 3653 2694 3691 2708
rect 3619 2660 3653 2674
rect 3687 2674 3691 2694
rect 3725 2674 3755 2708
rect 3687 2660 3755 2674
rect 3517 2628 3755 2660
rect 3517 2594 3547 2628
rect 3581 2594 3619 2628
rect 3653 2594 3691 2628
rect 3725 2594 3755 2628
rect 3517 2556 3755 2594
rect 3517 2540 3619 2556
rect 3653 2540 3755 2556
rect 3551 2518 3619 2540
rect 3653 2518 3721 2540
rect 3517 2472 3547 2506
rect 3725 2472 3755 2506
rect 3517 2404 3547 2438
rect 3725 2404 3755 2438
rect 3517 2336 3547 2370
rect 3725 2336 3755 2370
rect 3517 2268 3547 2302
rect 3725 2268 3755 2302
rect 3517 2200 3547 2234
rect 3725 2200 3755 2234
rect 3517 2132 3547 2166
rect 3725 2132 3755 2166
rect 3517 2064 3547 2098
rect 3725 2064 3755 2098
rect 3517 1996 3547 2030
rect 3725 1996 3755 2030
rect 3517 1928 3547 1962
rect 3725 1928 3755 1962
rect 3517 1860 3547 1894
rect 3725 1860 3755 1894
rect 3517 1792 3547 1826
rect 3725 1792 3755 1826
rect 3517 1724 3547 1758
rect 3725 1724 3755 1758
rect 3517 1656 3547 1690
rect 3725 1656 3755 1690
rect 3517 1620 3547 1622
rect 3725 1620 3755 1622
rect 3517 1586 3619 1620
rect 3653 1586 3755 1620
rect 3517 1536 3755 1586
rect 3857 3104 3977 4200
rect 4287 4308 4407 4324
rect 4287 4274 4330 4308
rect 4364 4274 4407 4308
rect 4287 4234 4407 4274
rect 4287 4200 4330 4234
rect 4364 4200 4407 4234
rect 3857 3070 3900 3104
rect 3934 3070 3977 3104
rect 3857 3026 3977 3070
rect 3857 2992 3900 3026
rect 3934 2992 3977 3026
rect 3857 2948 3977 2992
rect 3857 2914 3900 2948
rect 3934 2914 3977 2948
rect 3857 2870 3977 2914
rect 3857 2836 3900 2870
rect 3934 2836 3977 2870
rect 3857 2792 3977 2836
rect 3857 2758 3900 2792
rect 3934 2758 3977 2792
rect 3857 2713 3977 2758
rect 3857 2679 3900 2713
rect 3934 2679 3977 2713
rect 3857 2634 3977 2679
rect 3857 2600 3900 2634
rect 3934 2600 3977 2634
rect 3295 1470 3338 1504
rect 3372 1470 3415 1504
rect 3295 1430 3415 1470
rect 3295 1396 3338 1430
rect 3372 1396 3415 1430
rect 3295 1250 3415 1396
rect 3295 1144 3302 1250
rect 3408 1144 3415 1250
rect 3857 1504 3977 2600
rect 4042 4064 4043 4098
rect 4077 4082 4115 4098
rect 4077 4064 4079 4082
rect 4042 4048 4079 4064
rect 4113 4064 4115 4082
rect 4149 4082 4187 4098
rect 4149 4064 4151 4082
rect 4113 4048 4151 4064
rect 4185 4064 4187 4082
rect 4221 4064 4222 4098
rect 4185 4048 4222 4064
rect 4042 4025 4222 4048
rect 4042 3991 4043 4025
rect 4077 4014 4115 4025
rect 4077 3991 4079 4014
rect 4042 3980 4079 3991
rect 4113 3991 4115 4014
rect 4149 4014 4187 4025
rect 4149 3991 4151 4014
rect 4113 3980 4151 3991
rect 4185 3991 4187 4014
rect 4221 3991 4222 4025
rect 4185 3980 4222 3991
rect 4042 3952 4222 3980
rect 4042 3918 4043 3952
rect 4077 3946 4115 3952
rect 4077 3918 4079 3946
rect 4042 3912 4079 3918
rect 4113 3918 4115 3946
rect 4149 3946 4187 3952
rect 4149 3918 4151 3946
rect 4113 3912 4151 3918
rect 4185 3918 4187 3946
rect 4221 3918 4222 3952
rect 4185 3912 4222 3918
rect 4042 3879 4222 3912
rect 4042 3845 4043 3879
rect 4077 3878 4115 3879
rect 4077 3845 4079 3878
rect 4042 3844 4079 3845
rect 4113 3845 4115 3878
rect 4149 3878 4187 3879
rect 4149 3845 4151 3878
rect 4113 3844 4151 3845
rect 4185 3845 4187 3878
rect 4221 3845 4222 3879
rect 4185 3844 4222 3845
rect 4042 3810 4222 3844
rect 4042 3806 4079 3810
rect 4042 3772 4043 3806
rect 4077 3776 4079 3806
rect 4113 3806 4151 3810
rect 4113 3776 4115 3806
rect 4077 3772 4115 3776
rect 4149 3776 4151 3806
rect 4185 3806 4222 3810
rect 4185 3776 4187 3806
rect 4149 3772 4187 3776
rect 4221 3772 4222 3806
rect 4042 3742 4222 3772
rect 4042 3733 4079 3742
rect 4042 3699 4043 3733
rect 4077 3708 4079 3733
rect 4113 3733 4151 3742
rect 4113 3708 4115 3733
rect 4077 3699 4115 3708
rect 4149 3708 4151 3733
rect 4185 3733 4222 3742
rect 4185 3708 4187 3733
rect 4149 3699 4187 3708
rect 4221 3699 4222 3733
rect 4042 3674 4222 3699
rect 4042 3660 4079 3674
rect 4042 3626 4043 3660
rect 4077 3640 4079 3660
rect 4113 3660 4151 3674
rect 4113 3640 4115 3660
rect 4077 3626 4115 3640
rect 4149 3640 4151 3660
rect 4185 3660 4222 3674
rect 4185 3640 4187 3660
rect 4149 3626 4187 3640
rect 4221 3626 4222 3660
rect 4042 3606 4222 3626
rect 4042 3587 4079 3606
rect 4042 3553 4043 3587
rect 4077 3572 4079 3587
rect 4113 3587 4151 3606
rect 4113 3572 4115 3587
rect 4077 3553 4115 3572
rect 4149 3572 4151 3587
rect 4185 3587 4222 3606
rect 4185 3572 4187 3587
rect 4149 3553 4187 3572
rect 4221 3553 4222 3587
rect 4042 3538 4222 3553
rect 4042 3514 4079 3538
rect 4042 3480 4043 3514
rect 4077 3504 4079 3514
rect 4113 3514 4151 3538
rect 4113 3504 4115 3514
rect 4077 3480 4115 3504
rect 4149 3504 4151 3514
rect 4185 3514 4222 3538
rect 4185 3504 4187 3514
rect 4149 3480 4187 3504
rect 4221 3480 4222 3514
rect 4042 3470 4222 3480
rect 4042 3441 4079 3470
rect 4042 3407 4043 3441
rect 4077 3436 4079 3441
rect 4113 3441 4151 3470
rect 4113 3436 4115 3441
rect 4077 3407 4115 3436
rect 4149 3436 4151 3441
rect 4185 3441 4222 3470
rect 4185 3436 4187 3441
rect 4149 3407 4187 3436
rect 4221 3407 4222 3441
rect 4042 3402 4222 3407
rect 4042 3368 4079 3402
rect 4113 3368 4151 3402
rect 4185 3368 4222 3402
rect 4042 3334 4043 3368
rect 4077 3334 4115 3368
rect 4149 3334 4187 3368
rect 4221 3334 4222 3368
rect 4042 3300 4079 3334
rect 4113 3300 4151 3334
rect 4185 3300 4222 3334
rect 4042 3295 4222 3300
rect 4042 3261 4043 3295
rect 4077 3266 4115 3295
rect 4077 3261 4079 3266
rect 4042 3232 4079 3261
rect 4113 3261 4115 3266
rect 4149 3266 4187 3295
rect 4149 3261 4151 3266
rect 4113 3232 4151 3261
rect 4185 3261 4187 3266
rect 4221 3261 4222 3295
rect 4185 3232 4222 3261
rect 4042 3222 4222 3232
rect 4042 3188 4043 3222
rect 4077 3198 4115 3222
rect 4077 3188 4079 3198
rect 4042 3164 4079 3188
rect 4113 3188 4115 3198
rect 4149 3198 4187 3222
rect 4149 3188 4151 3198
rect 4113 3164 4151 3188
rect 4185 3188 4187 3198
rect 4221 3188 4222 3222
rect 4185 3164 4222 3188
rect 4042 3149 4222 3164
rect 4042 3115 4043 3149
rect 4077 3115 4115 3149
rect 4149 3115 4187 3149
rect 4221 3115 4222 3149
rect 4042 3076 4222 3115
rect 4042 3042 4043 3076
rect 4077 3042 4115 3076
rect 4149 3042 4187 3076
rect 4221 3042 4222 3076
rect 4042 3003 4222 3042
rect 4042 2969 4043 3003
rect 4077 2969 4115 3003
rect 4149 2969 4187 3003
rect 4221 2969 4222 3003
rect 4042 2930 4222 2969
rect 4042 2896 4043 2930
rect 4077 2896 4115 2930
rect 4149 2896 4187 2930
rect 4221 2896 4222 2930
rect 4042 2857 4222 2896
rect 4042 2823 4043 2857
rect 4077 2823 4115 2857
rect 4149 2823 4187 2857
rect 4221 2823 4222 2857
rect 4042 2784 4222 2823
rect 4042 2750 4043 2784
rect 4077 2750 4115 2784
rect 4149 2750 4187 2784
rect 4221 2750 4222 2784
rect 4042 2711 4222 2750
rect 4042 2677 4043 2711
rect 4077 2677 4115 2711
rect 4149 2677 4187 2711
rect 4221 2677 4222 2711
rect 4042 2638 4222 2677
rect 4042 2604 4043 2638
rect 4077 2604 4115 2638
rect 4149 2604 4187 2638
rect 4221 2604 4222 2638
rect 4042 2565 4222 2604
rect 4042 2531 4043 2565
rect 4077 2531 4115 2565
rect 4149 2531 4187 2565
rect 4221 2531 4222 2565
rect 4042 2492 4222 2531
rect 4042 2458 4043 2492
rect 4077 2482 4115 2492
rect 4077 2458 4079 2482
rect 4042 2448 4079 2458
rect 4113 2458 4115 2482
rect 4149 2482 4187 2492
rect 4149 2458 4151 2482
rect 4113 2448 4151 2458
rect 4185 2458 4187 2482
rect 4221 2458 4222 2492
rect 4185 2448 4222 2458
rect 4042 2419 4222 2448
rect 4042 2385 4043 2419
rect 4077 2414 4115 2419
rect 4077 2385 4079 2414
rect 4042 2380 4079 2385
rect 4113 2385 4115 2414
rect 4149 2414 4187 2419
rect 4149 2385 4151 2414
rect 4113 2380 4151 2385
rect 4185 2385 4187 2414
rect 4221 2385 4222 2419
rect 4185 2380 4222 2385
rect 4042 2346 4222 2380
rect 4042 2312 4043 2346
rect 4077 2312 4079 2346
rect 4113 2312 4115 2346
rect 4149 2312 4151 2346
rect 4185 2312 4187 2346
rect 4221 2312 4222 2346
rect 4042 2278 4222 2312
rect 4042 2273 4079 2278
rect 4042 2239 4043 2273
rect 4077 2244 4079 2273
rect 4113 2273 4151 2278
rect 4113 2244 4115 2273
rect 4077 2239 4115 2244
rect 4149 2244 4151 2273
rect 4185 2273 4222 2278
rect 4185 2244 4187 2273
rect 4149 2239 4187 2244
rect 4221 2239 4222 2273
rect 4042 2210 4222 2239
rect 4042 2200 4079 2210
rect 4042 2166 4043 2200
rect 4077 2176 4079 2200
rect 4113 2200 4151 2210
rect 4113 2176 4115 2200
rect 4077 2166 4115 2176
rect 4149 2176 4151 2200
rect 4185 2200 4222 2210
rect 4185 2176 4187 2200
rect 4149 2166 4187 2176
rect 4221 2166 4222 2200
rect 4042 2142 4222 2166
rect 4042 2126 4079 2142
rect 4042 2092 4043 2126
rect 4077 2108 4079 2126
rect 4113 2126 4151 2142
rect 4113 2108 4115 2126
rect 4077 2092 4115 2108
rect 4149 2108 4151 2126
rect 4185 2126 4222 2142
rect 4185 2108 4187 2126
rect 4149 2092 4187 2108
rect 4221 2092 4222 2126
rect 4042 2074 4222 2092
rect 4042 2052 4079 2074
rect 4042 2018 4043 2052
rect 4077 2040 4079 2052
rect 4113 2052 4151 2074
rect 4113 2040 4115 2052
rect 4077 2018 4115 2040
rect 4149 2040 4151 2052
rect 4185 2052 4222 2074
rect 4185 2040 4187 2052
rect 4149 2018 4187 2040
rect 4221 2018 4222 2052
rect 4042 2006 4222 2018
rect 4042 1978 4079 2006
rect 4042 1944 4043 1978
rect 4077 1972 4079 1978
rect 4113 1978 4151 2006
rect 4113 1972 4115 1978
rect 4077 1944 4115 1972
rect 4149 1972 4151 1978
rect 4185 1978 4222 2006
rect 4185 1972 4187 1978
rect 4149 1944 4187 1972
rect 4221 1944 4222 1978
rect 4042 1938 4222 1944
rect 4042 1904 4079 1938
rect 4113 1904 4151 1938
rect 4185 1904 4222 1938
rect 4042 1870 4043 1904
rect 4077 1870 4115 1904
rect 4149 1870 4187 1904
rect 4221 1870 4222 1904
rect 4042 1836 4079 1870
rect 4113 1836 4151 1870
rect 4185 1836 4222 1870
rect 4042 1830 4222 1836
rect 4042 1796 4043 1830
rect 4077 1802 4115 1830
rect 4077 1796 4079 1802
rect 4042 1768 4079 1796
rect 4113 1796 4115 1802
rect 4149 1802 4187 1830
rect 4149 1796 4151 1802
rect 4113 1768 4151 1796
rect 4185 1796 4187 1802
rect 4221 1796 4222 1830
rect 4185 1768 4222 1796
rect 4042 1756 4222 1768
rect 4042 1722 4043 1756
rect 4077 1734 4115 1756
rect 4077 1722 4079 1734
rect 4042 1700 4079 1722
rect 4113 1722 4115 1734
rect 4149 1734 4187 1756
rect 4149 1722 4151 1734
rect 4113 1700 4151 1722
rect 4185 1722 4187 1734
rect 4221 1722 4222 1756
rect 4185 1700 4222 1722
rect 4042 1682 4222 1700
rect 4042 1648 4043 1682
rect 4077 1666 4115 1682
rect 4077 1648 4079 1666
rect 4042 1632 4079 1648
rect 4113 1648 4115 1666
rect 4149 1666 4187 1682
rect 4149 1648 4151 1666
rect 4113 1632 4151 1648
rect 4185 1648 4187 1666
rect 4221 1648 4222 1682
rect 4185 1632 4222 1648
rect 4042 1608 4222 1632
rect 4042 1574 4043 1608
rect 4077 1598 4115 1608
rect 4077 1574 4079 1598
rect 4042 1564 4079 1574
rect 4113 1574 4115 1598
rect 4149 1598 4187 1608
rect 4149 1574 4151 1598
rect 4113 1564 4151 1574
rect 4185 1574 4187 1598
rect 4221 1574 4222 1608
rect 4185 1564 4222 1574
rect 4042 1548 4222 1564
rect 4287 3104 4407 4200
rect 4849 4308 4969 4324
rect 4849 4274 4892 4308
rect 4926 4274 4969 4308
rect 4849 4234 4969 4274
rect 4849 4200 4892 4234
rect 4926 4200 4969 4234
rect 4287 3070 4330 3104
rect 4364 3070 4407 3104
rect 4287 3026 4407 3070
rect 4287 2992 4330 3026
rect 4364 2992 4407 3026
rect 4287 2948 4407 2992
rect 4287 2914 4330 2948
rect 4364 2914 4407 2948
rect 4287 2870 4407 2914
rect 4287 2836 4330 2870
rect 4364 2836 4407 2870
rect 4287 2792 4407 2836
rect 4287 2758 4330 2792
rect 4364 2758 4407 2792
rect 4287 2713 4407 2758
rect 4287 2679 4330 2713
rect 4364 2679 4407 2713
rect 4287 2634 4407 2679
rect 4287 2600 4330 2634
rect 4364 2600 4407 2634
rect 3857 1470 3900 1504
rect 3934 1470 3977 1504
rect 3857 1430 3977 1470
rect 3857 1396 3900 1430
rect 3934 1396 3977 1430
rect 3857 1250 3977 1396
rect 3857 1144 3864 1250
rect 3970 1144 3977 1250
rect 4287 1504 4407 2600
rect 4509 4092 4611 4118
rect 4645 4092 4747 4118
rect 4509 4082 4539 4092
rect 4717 4082 4747 4092
rect 4509 4014 4539 4048
rect 4717 4014 4747 4048
rect 4509 3946 4539 3980
rect 4717 3946 4747 3980
rect 4509 3878 4539 3912
rect 4717 3878 4747 3912
rect 4509 3810 4539 3844
rect 4717 3810 4747 3844
rect 4509 3742 4539 3776
rect 4717 3742 4747 3776
rect 4509 3674 4539 3708
rect 4717 3674 4747 3708
rect 4509 3606 4539 3640
rect 4717 3606 4747 3640
rect 4509 3538 4539 3572
rect 4717 3538 4747 3572
rect 4509 3470 4539 3504
rect 4717 3470 4747 3504
rect 4509 3402 4539 3436
rect 4717 3402 4747 3436
rect 4509 3334 4539 3368
rect 4717 3334 4747 3368
rect 4509 3266 4539 3300
rect 4717 3266 4747 3300
rect 4509 3198 4539 3232
rect 4717 3198 4747 3232
rect 4543 3164 4611 3194
rect 4645 3164 4713 3194
rect 4509 3148 4611 3164
rect 4645 3148 4747 3164
rect 4509 3108 4747 3148
rect 4509 3074 4539 3108
rect 4573 3074 4611 3108
rect 4645 3074 4683 3108
rect 4717 3074 4747 3108
rect 4509 3044 4747 3074
rect 4509 3028 4577 3044
rect 4509 2994 4539 3028
rect 4573 3010 4577 3028
rect 4611 3028 4645 3044
rect 4573 2994 4611 3010
rect 4679 3028 4747 3044
rect 4679 3010 4683 3028
rect 4645 2994 4683 3010
rect 4717 2994 4747 3028
rect 4509 2974 4747 2994
rect 4509 2948 4577 2974
rect 4509 2914 4539 2948
rect 4573 2940 4577 2948
rect 4611 2948 4645 2974
rect 4573 2914 4611 2940
rect 4679 2948 4747 2974
rect 4679 2940 4683 2948
rect 4645 2914 4683 2940
rect 4717 2914 4747 2948
rect 4509 2904 4747 2914
rect 4509 2870 4577 2904
rect 4611 2870 4645 2904
rect 4679 2870 4747 2904
rect 4509 2868 4747 2870
rect 4509 2834 4539 2868
rect 4573 2834 4611 2868
rect 4645 2834 4683 2868
rect 4717 2834 4747 2868
rect 4509 2800 4577 2834
rect 4611 2800 4645 2834
rect 4679 2800 4747 2834
rect 4509 2788 4747 2800
rect 4509 2754 4539 2788
rect 4573 2764 4611 2788
rect 4573 2754 4577 2764
rect 4509 2730 4577 2754
rect 4645 2764 4683 2788
rect 4611 2730 4645 2754
rect 4679 2754 4683 2764
rect 4717 2754 4747 2788
rect 4679 2730 4747 2754
rect 4509 2708 4747 2730
rect 4509 2674 4539 2708
rect 4573 2694 4611 2708
rect 4573 2674 4577 2694
rect 4509 2660 4577 2674
rect 4645 2694 4683 2708
rect 4611 2660 4645 2674
rect 4679 2674 4683 2694
rect 4717 2674 4747 2708
rect 4679 2660 4747 2674
rect 4509 2628 4747 2660
rect 4509 2594 4539 2628
rect 4573 2594 4611 2628
rect 4645 2594 4683 2628
rect 4717 2594 4747 2628
rect 4509 2556 4747 2594
rect 4509 2540 4611 2556
rect 4645 2540 4747 2556
rect 4543 2518 4611 2540
rect 4645 2518 4713 2540
rect 4509 2472 4539 2506
rect 4717 2472 4747 2506
rect 4509 2404 4539 2438
rect 4717 2404 4747 2438
rect 4509 2336 4539 2370
rect 4717 2336 4747 2370
rect 4509 2268 4539 2302
rect 4717 2268 4747 2302
rect 4509 2200 4539 2234
rect 4717 2200 4747 2234
rect 4509 2132 4539 2166
rect 4717 2132 4747 2166
rect 4509 2064 4539 2098
rect 4717 2064 4747 2098
rect 4509 1996 4539 2030
rect 4717 1996 4747 2030
rect 4509 1928 4539 1962
rect 4717 1928 4747 1962
rect 4509 1860 4539 1894
rect 4717 1860 4747 1894
rect 4509 1792 4539 1826
rect 4717 1792 4747 1826
rect 4509 1724 4539 1758
rect 4717 1724 4747 1758
rect 4509 1656 4539 1690
rect 4717 1656 4747 1690
rect 4509 1620 4539 1622
rect 4717 1620 4747 1622
rect 4509 1586 4611 1620
rect 4645 1586 4747 1620
rect 4509 1536 4747 1586
rect 4849 3104 4969 4200
rect 5279 4308 5399 4324
rect 5279 4274 5322 4308
rect 5356 4274 5399 4308
rect 5279 4234 5399 4274
rect 5279 4200 5322 4234
rect 5356 4200 5399 4234
rect 4849 3070 4892 3104
rect 4926 3070 4969 3104
rect 4849 3026 4969 3070
rect 4849 2992 4892 3026
rect 4926 2992 4969 3026
rect 4849 2948 4969 2992
rect 4849 2914 4892 2948
rect 4926 2914 4969 2948
rect 4849 2870 4969 2914
rect 4849 2836 4892 2870
rect 4926 2836 4969 2870
rect 4849 2792 4969 2836
rect 4849 2758 4892 2792
rect 4926 2758 4969 2792
rect 4849 2713 4969 2758
rect 4849 2679 4892 2713
rect 4926 2679 4969 2713
rect 4849 2634 4969 2679
rect 4849 2600 4892 2634
rect 4926 2600 4969 2634
rect 4287 1470 4330 1504
rect 4364 1470 4407 1504
rect 4287 1430 4407 1470
rect 4287 1396 4330 1430
rect 4364 1396 4407 1430
rect 4287 1250 4407 1396
rect 4287 1144 4294 1250
rect 4400 1144 4407 1250
rect 4849 1504 4969 2600
rect 5034 4064 5035 4098
rect 5069 4082 5107 4098
rect 5069 4064 5071 4082
rect 5034 4048 5071 4064
rect 5105 4064 5107 4082
rect 5141 4082 5179 4098
rect 5141 4064 5143 4082
rect 5105 4048 5143 4064
rect 5177 4064 5179 4082
rect 5213 4064 5214 4098
rect 5177 4048 5214 4064
rect 5034 4025 5214 4048
rect 5034 3991 5035 4025
rect 5069 4014 5107 4025
rect 5069 3991 5071 4014
rect 5034 3980 5071 3991
rect 5105 3991 5107 4014
rect 5141 4014 5179 4025
rect 5141 3991 5143 4014
rect 5105 3980 5143 3991
rect 5177 3991 5179 4014
rect 5213 3991 5214 4025
rect 5177 3980 5214 3991
rect 5034 3952 5214 3980
rect 5034 3918 5035 3952
rect 5069 3946 5107 3952
rect 5069 3918 5071 3946
rect 5034 3912 5071 3918
rect 5105 3918 5107 3946
rect 5141 3946 5179 3952
rect 5141 3918 5143 3946
rect 5105 3912 5143 3918
rect 5177 3918 5179 3946
rect 5213 3918 5214 3952
rect 5177 3912 5214 3918
rect 5034 3879 5214 3912
rect 5034 3845 5035 3879
rect 5069 3878 5107 3879
rect 5069 3845 5071 3878
rect 5034 3844 5071 3845
rect 5105 3845 5107 3878
rect 5141 3878 5179 3879
rect 5141 3845 5143 3878
rect 5105 3844 5143 3845
rect 5177 3845 5179 3878
rect 5213 3845 5214 3879
rect 5177 3844 5214 3845
rect 5034 3810 5214 3844
rect 5034 3806 5071 3810
rect 5034 3772 5035 3806
rect 5069 3776 5071 3806
rect 5105 3806 5143 3810
rect 5105 3776 5107 3806
rect 5069 3772 5107 3776
rect 5141 3776 5143 3806
rect 5177 3806 5214 3810
rect 5177 3776 5179 3806
rect 5141 3772 5179 3776
rect 5213 3772 5214 3806
rect 5034 3742 5214 3772
rect 5034 3733 5071 3742
rect 5034 3699 5035 3733
rect 5069 3708 5071 3733
rect 5105 3733 5143 3742
rect 5105 3708 5107 3733
rect 5069 3699 5107 3708
rect 5141 3708 5143 3733
rect 5177 3733 5214 3742
rect 5177 3708 5179 3733
rect 5141 3699 5179 3708
rect 5213 3699 5214 3733
rect 5034 3674 5214 3699
rect 5034 3660 5071 3674
rect 5034 3626 5035 3660
rect 5069 3640 5071 3660
rect 5105 3660 5143 3674
rect 5105 3640 5107 3660
rect 5069 3626 5107 3640
rect 5141 3640 5143 3660
rect 5177 3660 5214 3674
rect 5177 3640 5179 3660
rect 5141 3626 5179 3640
rect 5213 3626 5214 3660
rect 5034 3606 5214 3626
rect 5034 3587 5071 3606
rect 5034 3553 5035 3587
rect 5069 3572 5071 3587
rect 5105 3587 5143 3606
rect 5105 3572 5107 3587
rect 5069 3553 5107 3572
rect 5141 3572 5143 3587
rect 5177 3587 5214 3606
rect 5177 3572 5179 3587
rect 5141 3553 5179 3572
rect 5213 3553 5214 3587
rect 5034 3538 5214 3553
rect 5034 3514 5071 3538
rect 5034 3480 5035 3514
rect 5069 3504 5071 3514
rect 5105 3514 5143 3538
rect 5105 3504 5107 3514
rect 5069 3480 5107 3504
rect 5141 3504 5143 3514
rect 5177 3514 5214 3538
rect 5177 3504 5179 3514
rect 5141 3480 5179 3504
rect 5213 3480 5214 3514
rect 5034 3470 5214 3480
rect 5034 3441 5071 3470
rect 5034 3407 5035 3441
rect 5069 3436 5071 3441
rect 5105 3441 5143 3470
rect 5105 3436 5107 3441
rect 5069 3407 5107 3436
rect 5141 3436 5143 3441
rect 5177 3441 5214 3470
rect 5177 3436 5179 3441
rect 5141 3407 5179 3436
rect 5213 3407 5214 3441
rect 5034 3402 5214 3407
rect 5034 3368 5071 3402
rect 5105 3368 5143 3402
rect 5177 3368 5214 3402
rect 5034 3334 5035 3368
rect 5069 3334 5107 3368
rect 5141 3334 5179 3368
rect 5213 3334 5214 3368
rect 5034 3300 5071 3334
rect 5105 3300 5143 3334
rect 5177 3300 5214 3334
rect 5034 3295 5214 3300
rect 5034 3261 5035 3295
rect 5069 3266 5107 3295
rect 5069 3261 5071 3266
rect 5034 3232 5071 3261
rect 5105 3261 5107 3266
rect 5141 3266 5179 3295
rect 5141 3261 5143 3266
rect 5105 3232 5143 3261
rect 5177 3261 5179 3266
rect 5213 3261 5214 3295
rect 5177 3232 5214 3261
rect 5034 3222 5214 3232
rect 5034 3188 5035 3222
rect 5069 3198 5107 3222
rect 5069 3188 5071 3198
rect 5034 3164 5071 3188
rect 5105 3188 5107 3198
rect 5141 3198 5179 3222
rect 5141 3188 5143 3198
rect 5105 3164 5143 3188
rect 5177 3188 5179 3198
rect 5213 3188 5214 3222
rect 5177 3164 5214 3188
rect 5034 3149 5214 3164
rect 5034 3115 5035 3149
rect 5069 3115 5107 3149
rect 5141 3115 5179 3149
rect 5213 3115 5214 3149
rect 5034 3076 5214 3115
rect 5034 3042 5035 3076
rect 5069 3042 5107 3076
rect 5141 3042 5179 3076
rect 5213 3042 5214 3076
rect 5034 3003 5214 3042
rect 5034 2969 5035 3003
rect 5069 2969 5107 3003
rect 5141 2969 5179 3003
rect 5213 2969 5214 3003
rect 5034 2930 5214 2969
rect 5034 2896 5035 2930
rect 5069 2896 5107 2930
rect 5141 2896 5179 2930
rect 5213 2896 5214 2930
rect 5034 2857 5214 2896
rect 5034 2823 5035 2857
rect 5069 2823 5107 2857
rect 5141 2823 5179 2857
rect 5213 2823 5214 2857
rect 5034 2784 5214 2823
rect 5034 2750 5035 2784
rect 5069 2750 5107 2784
rect 5141 2750 5179 2784
rect 5213 2750 5214 2784
rect 5034 2711 5214 2750
rect 5034 2677 5035 2711
rect 5069 2677 5107 2711
rect 5141 2677 5179 2711
rect 5213 2677 5214 2711
rect 5034 2638 5214 2677
rect 5034 2604 5035 2638
rect 5069 2604 5107 2638
rect 5141 2604 5179 2638
rect 5213 2604 5214 2638
rect 5034 2565 5214 2604
rect 5034 2531 5035 2565
rect 5069 2531 5107 2565
rect 5141 2531 5179 2565
rect 5213 2531 5214 2565
rect 5034 2492 5214 2531
rect 5034 2458 5035 2492
rect 5069 2482 5107 2492
rect 5069 2458 5071 2482
rect 5034 2448 5071 2458
rect 5105 2458 5107 2482
rect 5141 2482 5179 2492
rect 5141 2458 5143 2482
rect 5105 2448 5143 2458
rect 5177 2458 5179 2482
rect 5213 2458 5214 2492
rect 5177 2448 5214 2458
rect 5034 2419 5214 2448
rect 5034 2385 5035 2419
rect 5069 2414 5107 2419
rect 5069 2385 5071 2414
rect 5034 2380 5071 2385
rect 5105 2385 5107 2414
rect 5141 2414 5179 2419
rect 5141 2385 5143 2414
rect 5105 2380 5143 2385
rect 5177 2385 5179 2414
rect 5213 2385 5214 2419
rect 5177 2380 5214 2385
rect 5034 2346 5214 2380
rect 5034 2312 5035 2346
rect 5069 2312 5071 2346
rect 5105 2312 5107 2346
rect 5141 2312 5143 2346
rect 5177 2312 5179 2346
rect 5213 2312 5214 2346
rect 5034 2278 5214 2312
rect 5034 2273 5071 2278
rect 5034 2239 5035 2273
rect 5069 2244 5071 2273
rect 5105 2273 5143 2278
rect 5105 2244 5107 2273
rect 5069 2239 5107 2244
rect 5141 2244 5143 2273
rect 5177 2273 5214 2278
rect 5177 2244 5179 2273
rect 5141 2239 5179 2244
rect 5213 2239 5214 2273
rect 5034 2210 5214 2239
rect 5034 2200 5071 2210
rect 5034 2166 5035 2200
rect 5069 2176 5071 2200
rect 5105 2200 5143 2210
rect 5105 2176 5107 2200
rect 5069 2166 5107 2176
rect 5141 2176 5143 2200
rect 5177 2200 5214 2210
rect 5177 2176 5179 2200
rect 5141 2166 5179 2176
rect 5213 2166 5214 2200
rect 5034 2142 5214 2166
rect 5034 2126 5071 2142
rect 5034 2092 5035 2126
rect 5069 2108 5071 2126
rect 5105 2126 5143 2142
rect 5105 2108 5107 2126
rect 5069 2092 5107 2108
rect 5141 2108 5143 2126
rect 5177 2126 5214 2142
rect 5177 2108 5179 2126
rect 5141 2092 5179 2108
rect 5213 2092 5214 2126
rect 5034 2074 5214 2092
rect 5034 2052 5071 2074
rect 5034 2018 5035 2052
rect 5069 2040 5071 2052
rect 5105 2052 5143 2074
rect 5105 2040 5107 2052
rect 5069 2018 5107 2040
rect 5141 2040 5143 2052
rect 5177 2052 5214 2074
rect 5177 2040 5179 2052
rect 5141 2018 5179 2040
rect 5213 2018 5214 2052
rect 5034 2006 5214 2018
rect 5034 1978 5071 2006
rect 5034 1944 5035 1978
rect 5069 1972 5071 1978
rect 5105 1978 5143 2006
rect 5105 1972 5107 1978
rect 5069 1944 5107 1972
rect 5141 1972 5143 1978
rect 5177 1978 5214 2006
rect 5177 1972 5179 1978
rect 5141 1944 5179 1972
rect 5213 1944 5214 1978
rect 5034 1938 5214 1944
rect 5034 1904 5071 1938
rect 5105 1904 5143 1938
rect 5177 1904 5214 1938
rect 5034 1870 5035 1904
rect 5069 1870 5107 1904
rect 5141 1870 5179 1904
rect 5213 1870 5214 1904
rect 5034 1836 5071 1870
rect 5105 1836 5143 1870
rect 5177 1836 5214 1870
rect 5034 1830 5214 1836
rect 5034 1796 5035 1830
rect 5069 1802 5107 1830
rect 5069 1796 5071 1802
rect 5034 1768 5071 1796
rect 5105 1796 5107 1802
rect 5141 1802 5179 1830
rect 5141 1796 5143 1802
rect 5105 1768 5143 1796
rect 5177 1796 5179 1802
rect 5213 1796 5214 1830
rect 5177 1768 5214 1796
rect 5034 1756 5214 1768
rect 5034 1722 5035 1756
rect 5069 1734 5107 1756
rect 5069 1722 5071 1734
rect 5034 1700 5071 1722
rect 5105 1722 5107 1734
rect 5141 1734 5179 1756
rect 5141 1722 5143 1734
rect 5105 1700 5143 1722
rect 5177 1722 5179 1734
rect 5213 1722 5214 1756
rect 5177 1700 5214 1722
rect 5034 1682 5214 1700
rect 5034 1648 5035 1682
rect 5069 1666 5107 1682
rect 5069 1648 5071 1666
rect 5034 1632 5071 1648
rect 5105 1648 5107 1666
rect 5141 1666 5179 1682
rect 5141 1648 5143 1666
rect 5105 1632 5143 1648
rect 5177 1648 5179 1666
rect 5213 1648 5214 1682
rect 5177 1632 5214 1648
rect 5034 1608 5214 1632
rect 5034 1574 5035 1608
rect 5069 1598 5107 1608
rect 5069 1574 5071 1598
rect 5034 1564 5071 1574
rect 5105 1574 5107 1598
rect 5141 1598 5179 1608
rect 5141 1574 5143 1598
rect 5105 1564 5143 1574
rect 5177 1574 5179 1598
rect 5213 1574 5214 1608
rect 5177 1564 5214 1574
rect 5034 1548 5214 1564
rect 5279 3104 5399 4200
rect 5841 4308 5961 4324
rect 5841 4274 5884 4308
rect 5918 4274 5961 4308
rect 5841 4234 5961 4274
rect 5841 4200 5884 4234
rect 5918 4200 5961 4234
rect 5279 3070 5322 3104
rect 5356 3070 5399 3104
rect 5279 3026 5399 3070
rect 5279 2992 5322 3026
rect 5356 2992 5399 3026
rect 5279 2948 5399 2992
rect 5279 2914 5322 2948
rect 5356 2914 5399 2948
rect 5279 2870 5399 2914
rect 5279 2836 5322 2870
rect 5356 2836 5399 2870
rect 5279 2792 5399 2836
rect 5279 2758 5322 2792
rect 5356 2758 5399 2792
rect 5279 2713 5399 2758
rect 5279 2679 5322 2713
rect 5356 2679 5399 2713
rect 5279 2634 5399 2679
rect 5279 2600 5322 2634
rect 5356 2600 5399 2634
rect 4849 1470 4892 1504
rect 4926 1470 4969 1504
rect 4849 1430 4969 1470
rect 4849 1396 4892 1430
rect 4926 1396 4969 1430
rect 4849 1250 4969 1396
rect 4849 1144 4856 1250
rect 4962 1144 4969 1250
rect 5279 1504 5399 2600
rect 5501 4092 5603 4118
rect 5637 4092 5739 4118
rect 5501 4082 5531 4092
rect 5709 4082 5739 4092
rect 5501 4014 5531 4048
rect 5709 4014 5739 4048
rect 5501 3946 5531 3980
rect 5709 3946 5739 3980
rect 5501 3878 5531 3912
rect 5709 3878 5739 3912
rect 5501 3810 5531 3844
rect 5709 3810 5739 3844
rect 5501 3742 5531 3776
rect 5709 3742 5739 3776
rect 5501 3674 5531 3708
rect 5709 3674 5739 3708
rect 5501 3606 5531 3640
rect 5709 3606 5739 3640
rect 5501 3538 5531 3572
rect 5709 3538 5739 3572
rect 5501 3470 5531 3504
rect 5709 3470 5739 3504
rect 5501 3402 5531 3436
rect 5709 3402 5739 3436
rect 5501 3334 5531 3368
rect 5709 3334 5739 3368
rect 5501 3266 5531 3300
rect 5709 3266 5739 3300
rect 5501 3198 5531 3232
rect 5709 3198 5739 3232
rect 5535 3164 5603 3194
rect 5637 3164 5705 3194
rect 5501 3148 5603 3164
rect 5637 3148 5739 3164
rect 5501 3108 5739 3148
rect 5501 3074 5531 3108
rect 5565 3074 5603 3108
rect 5637 3074 5675 3108
rect 5709 3074 5739 3108
rect 5501 3044 5739 3074
rect 5501 3028 5569 3044
rect 5501 2994 5531 3028
rect 5565 3010 5569 3028
rect 5603 3028 5637 3044
rect 5565 2994 5603 3010
rect 5671 3028 5739 3044
rect 5671 3010 5675 3028
rect 5637 2994 5675 3010
rect 5709 2994 5739 3028
rect 5501 2974 5739 2994
rect 5501 2948 5569 2974
rect 5501 2914 5531 2948
rect 5565 2940 5569 2948
rect 5603 2948 5637 2974
rect 5565 2914 5603 2940
rect 5671 2948 5739 2974
rect 5671 2940 5675 2948
rect 5637 2914 5675 2940
rect 5709 2914 5739 2948
rect 5501 2904 5739 2914
rect 5501 2870 5569 2904
rect 5603 2870 5637 2904
rect 5671 2870 5739 2904
rect 5501 2868 5739 2870
rect 5501 2834 5531 2868
rect 5565 2834 5603 2868
rect 5637 2834 5675 2868
rect 5709 2834 5739 2868
rect 5501 2800 5569 2834
rect 5603 2800 5637 2834
rect 5671 2800 5739 2834
rect 5501 2788 5739 2800
rect 5501 2754 5531 2788
rect 5565 2764 5603 2788
rect 5565 2754 5569 2764
rect 5501 2730 5569 2754
rect 5637 2764 5675 2788
rect 5603 2730 5637 2754
rect 5671 2754 5675 2764
rect 5709 2754 5739 2788
rect 5671 2730 5739 2754
rect 5501 2708 5739 2730
rect 5501 2674 5531 2708
rect 5565 2694 5603 2708
rect 5565 2674 5569 2694
rect 5501 2660 5569 2674
rect 5637 2694 5675 2708
rect 5603 2660 5637 2674
rect 5671 2674 5675 2694
rect 5709 2674 5739 2708
rect 5671 2660 5739 2674
rect 5501 2628 5739 2660
rect 5501 2594 5531 2628
rect 5565 2594 5603 2628
rect 5637 2594 5675 2628
rect 5709 2594 5739 2628
rect 5501 2556 5739 2594
rect 5501 2540 5603 2556
rect 5637 2540 5739 2556
rect 5535 2518 5603 2540
rect 5637 2518 5705 2540
rect 5501 2472 5531 2506
rect 5709 2472 5739 2506
rect 5501 2404 5531 2438
rect 5709 2404 5739 2438
rect 5501 2336 5531 2370
rect 5709 2336 5739 2370
rect 5501 2268 5531 2302
rect 5709 2268 5739 2302
rect 5501 2200 5531 2234
rect 5709 2200 5739 2234
rect 5501 2132 5531 2166
rect 5709 2132 5739 2166
rect 5501 2064 5531 2098
rect 5709 2064 5739 2098
rect 5501 1996 5531 2030
rect 5709 1996 5739 2030
rect 5501 1928 5531 1962
rect 5709 1928 5739 1962
rect 5501 1860 5531 1894
rect 5709 1860 5739 1894
rect 5501 1792 5531 1826
rect 5709 1792 5739 1826
rect 5501 1724 5531 1758
rect 5709 1724 5739 1758
rect 5501 1656 5531 1690
rect 5709 1656 5739 1690
rect 5501 1620 5531 1622
rect 5709 1620 5739 1622
rect 5501 1586 5603 1620
rect 5637 1586 5739 1620
rect 5501 1536 5739 1586
rect 5841 3104 5961 4200
rect 6271 4308 6391 4324
rect 6271 4274 6314 4308
rect 6348 4274 6391 4308
rect 6271 4234 6391 4274
rect 6271 4200 6314 4234
rect 6348 4200 6391 4234
rect 5841 3070 5884 3104
rect 5918 3070 5961 3104
rect 5841 3026 5961 3070
rect 5841 2992 5884 3026
rect 5918 2992 5961 3026
rect 5841 2948 5961 2992
rect 5841 2914 5884 2948
rect 5918 2914 5961 2948
rect 5841 2870 5961 2914
rect 5841 2836 5884 2870
rect 5918 2836 5961 2870
rect 5841 2792 5961 2836
rect 5841 2758 5884 2792
rect 5918 2758 5961 2792
rect 5841 2713 5961 2758
rect 5841 2679 5884 2713
rect 5918 2679 5961 2713
rect 5841 2634 5961 2679
rect 5841 2600 5884 2634
rect 5918 2600 5961 2634
rect 5279 1470 5322 1504
rect 5356 1470 5399 1504
rect 5279 1430 5399 1470
rect 5279 1396 5322 1430
rect 5356 1396 5399 1430
rect 5279 1250 5399 1396
rect 5279 1144 5286 1250
rect 5392 1144 5399 1250
rect 5841 1504 5961 2600
rect 6026 4064 6027 4098
rect 6061 4082 6099 4098
rect 6061 4064 6063 4082
rect 6026 4048 6063 4064
rect 6097 4064 6099 4082
rect 6133 4082 6171 4098
rect 6133 4064 6135 4082
rect 6097 4048 6135 4064
rect 6169 4064 6171 4082
rect 6205 4064 6206 4098
rect 6169 4048 6206 4064
rect 6026 4025 6206 4048
rect 6026 3991 6027 4025
rect 6061 4014 6099 4025
rect 6061 3991 6063 4014
rect 6026 3980 6063 3991
rect 6097 3991 6099 4014
rect 6133 4014 6171 4025
rect 6133 3991 6135 4014
rect 6097 3980 6135 3991
rect 6169 3991 6171 4014
rect 6205 3991 6206 4025
rect 6169 3980 6206 3991
rect 6026 3952 6206 3980
rect 6026 3918 6027 3952
rect 6061 3946 6099 3952
rect 6061 3918 6063 3946
rect 6026 3912 6063 3918
rect 6097 3918 6099 3946
rect 6133 3946 6171 3952
rect 6133 3918 6135 3946
rect 6097 3912 6135 3918
rect 6169 3918 6171 3946
rect 6205 3918 6206 3952
rect 6169 3912 6206 3918
rect 6026 3879 6206 3912
rect 6026 3845 6027 3879
rect 6061 3878 6099 3879
rect 6061 3845 6063 3878
rect 6026 3844 6063 3845
rect 6097 3845 6099 3878
rect 6133 3878 6171 3879
rect 6133 3845 6135 3878
rect 6097 3844 6135 3845
rect 6169 3845 6171 3878
rect 6205 3845 6206 3879
rect 6169 3844 6206 3845
rect 6026 3810 6206 3844
rect 6026 3806 6063 3810
rect 6026 3772 6027 3806
rect 6061 3776 6063 3806
rect 6097 3806 6135 3810
rect 6097 3776 6099 3806
rect 6061 3772 6099 3776
rect 6133 3776 6135 3806
rect 6169 3806 6206 3810
rect 6169 3776 6171 3806
rect 6133 3772 6171 3776
rect 6205 3772 6206 3806
rect 6026 3742 6206 3772
rect 6026 3733 6063 3742
rect 6026 3699 6027 3733
rect 6061 3708 6063 3733
rect 6097 3733 6135 3742
rect 6097 3708 6099 3733
rect 6061 3699 6099 3708
rect 6133 3708 6135 3733
rect 6169 3733 6206 3742
rect 6169 3708 6171 3733
rect 6133 3699 6171 3708
rect 6205 3699 6206 3733
rect 6026 3674 6206 3699
rect 6026 3660 6063 3674
rect 6026 3626 6027 3660
rect 6061 3640 6063 3660
rect 6097 3660 6135 3674
rect 6097 3640 6099 3660
rect 6061 3626 6099 3640
rect 6133 3640 6135 3660
rect 6169 3660 6206 3674
rect 6169 3640 6171 3660
rect 6133 3626 6171 3640
rect 6205 3626 6206 3660
rect 6026 3606 6206 3626
rect 6026 3587 6063 3606
rect 6026 3553 6027 3587
rect 6061 3572 6063 3587
rect 6097 3587 6135 3606
rect 6097 3572 6099 3587
rect 6061 3553 6099 3572
rect 6133 3572 6135 3587
rect 6169 3587 6206 3606
rect 6169 3572 6171 3587
rect 6133 3553 6171 3572
rect 6205 3553 6206 3587
rect 6026 3538 6206 3553
rect 6026 3514 6063 3538
rect 6026 3480 6027 3514
rect 6061 3504 6063 3514
rect 6097 3514 6135 3538
rect 6097 3504 6099 3514
rect 6061 3480 6099 3504
rect 6133 3504 6135 3514
rect 6169 3514 6206 3538
rect 6169 3504 6171 3514
rect 6133 3480 6171 3504
rect 6205 3480 6206 3514
rect 6026 3470 6206 3480
rect 6026 3441 6063 3470
rect 6026 3407 6027 3441
rect 6061 3436 6063 3441
rect 6097 3441 6135 3470
rect 6097 3436 6099 3441
rect 6061 3407 6099 3436
rect 6133 3436 6135 3441
rect 6169 3441 6206 3470
rect 6169 3436 6171 3441
rect 6133 3407 6171 3436
rect 6205 3407 6206 3441
rect 6026 3402 6206 3407
rect 6026 3368 6063 3402
rect 6097 3368 6135 3402
rect 6169 3368 6206 3402
rect 6026 3334 6027 3368
rect 6061 3334 6099 3368
rect 6133 3334 6171 3368
rect 6205 3334 6206 3368
rect 6026 3300 6063 3334
rect 6097 3300 6135 3334
rect 6169 3300 6206 3334
rect 6026 3295 6206 3300
rect 6026 3261 6027 3295
rect 6061 3266 6099 3295
rect 6061 3261 6063 3266
rect 6026 3232 6063 3261
rect 6097 3261 6099 3266
rect 6133 3266 6171 3295
rect 6133 3261 6135 3266
rect 6097 3232 6135 3261
rect 6169 3261 6171 3266
rect 6205 3261 6206 3295
rect 6169 3232 6206 3261
rect 6026 3222 6206 3232
rect 6026 3188 6027 3222
rect 6061 3198 6099 3222
rect 6061 3188 6063 3198
rect 6026 3164 6063 3188
rect 6097 3188 6099 3198
rect 6133 3198 6171 3222
rect 6133 3188 6135 3198
rect 6097 3164 6135 3188
rect 6169 3188 6171 3198
rect 6205 3188 6206 3222
rect 6169 3164 6206 3188
rect 6026 3149 6206 3164
rect 6026 3115 6027 3149
rect 6061 3115 6099 3149
rect 6133 3115 6171 3149
rect 6205 3115 6206 3149
rect 6026 3076 6206 3115
rect 6026 3042 6027 3076
rect 6061 3042 6099 3076
rect 6133 3042 6171 3076
rect 6205 3042 6206 3076
rect 6026 3003 6206 3042
rect 6026 2969 6027 3003
rect 6061 2969 6099 3003
rect 6133 2969 6171 3003
rect 6205 2969 6206 3003
rect 6026 2930 6206 2969
rect 6026 2896 6027 2930
rect 6061 2896 6099 2930
rect 6133 2896 6171 2930
rect 6205 2896 6206 2930
rect 6026 2857 6206 2896
rect 6026 2823 6027 2857
rect 6061 2823 6099 2857
rect 6133 2823 6171 2857
rect 6205 2823 6206 2857
rect 6026 2784 6206 2823
rect 6026 2750 6027 2784
rect 6061 2750 6099 2784
rect 6133 2750 6171 2784
rect 6205 2750 6206 2784
rect 6026 2711 6206 2750
rect 6026 2677 6027 2711
rect 6061 2677 6099 2711
rect 6133 2677 6171 2711
rect 6205 2677 6206 2711
rect 6026 2638 6206 2677
rect 6026 2604 6027 2638
rect 6061 2604 6099 2638
rect 6133 2604 6171 2638
rect 6205 2604 6206 2638
rect 6026 2565 6206 2604
rect 6026 2531 6027 2565
rect 6061 2531 6099 2565
rect 6133 2531 6171 2565
rect 6205 2531 6206 2565
rect 6026 2492 6206 2531
rect 6026 2458 6027 2492
rect 6061 2482 6099 2492
rect 6061 2458 6063 2482
rect 6026 2448 6063 2458
rect 6097 2458 6099 2482
rect 6133 2482 6171 2492
rect 6133 2458 6135 2482
rect 6097 2448 6135 2458
rect 6169 2458 6171 2482
rect 6205 2458 6206 2492
rect 6169 2448 6206 2458
rect 6026 2419 6206 2448
rect 6026 2385 6027 2419
rect 6061 2414 6099 2419
rect 6061 2385 6063 2414
rect 6026 2380 6063 2385
rect 6097 2385 6099 2414
rect 6133 2414 6171 2419
rect 6133 2385 6135 2414
rect 6097 2380 6135 2385
rect 6169 2385 6171 2414
rect 6205 2385 6206 2419
rect 6169 2380 6206 2385
rect 6026 2346 6206 2380
rect 6026 2312 6027 2346
rect 6061 2312 6063 2346
rect 6097 2312 6099 2346
rect 6133 2312 6135 2346
rect 6169 2312 6171 2346
rect 6205 2312 6206 2346
rect 6026 2278 6206 2312
rect 6026 2273 6063 2278
rect 6026 2239 6027 2273
rect 6061 2244 6063 2273
rect 6097 2273 6135 2278
rect 6097 2244 6099 2273
rect 6061 2239 6099 2244
rect 6133 2244 6135 2273
rect 6169 2273 6206 2278
rect 6169 2244 6171 2273
rect 6133 2239 6171 2244
rect 6205 2239 6206 2273
rect 6026 2210 6206 2239
rect 6026 2200 6063 2210
rect 6026 2166 6027 2200
rect 6061 2176 6063 2200
rect 6097 2200 6135 2210
rect 6097 2176 6099 2200
rect 6061 2166 6099 2176
rect 6133 2176 6135 2200
rect 6169 2200 6206 2210
rect 6169 2176 6171 2200
rect 6133 2166 6171 2176
rect 6205 2166 6206 2200
rect 6026 2142 6206 2166
rect 6026 2126 6063 2142
rect 6026 2092 6027 2126
rect 6061 2108 6063 2126
rect 6097 2126 6135 2142
rect 6097 2108 6099 2126
rect 6061 2092 6099 2108
rect 6133 2108 6135 2126
rect 6169 2126 6206 2142
rect 6169 2108 6171 2126
rect 6133 2092 6171 2108
rect 6205 2092 6206 2126
rect 6026 2074 6206 2092
rect 6026 2052 6063 2074
rect 6026 2018 6027 2052
rect 6061 2040 6063 2052
rect 6097 2052 6135 2074
rect 6097 2040 6099 2052
rect 6061 2018 6099 2040
rect 6133 2040 6135 2052
rect 6169 2052 6206 2074
rect 6169 2040 6171 2052
rect 6133 2018 6171 2040
rect 6205 2018 6206 2052
rect 6026 2006 6206 2018
rect 6026 1978 6063 2006
rect 6026 1944 6027 1978
rect 6061 1972 6063 1978
rect 6097 1978 6135 2006
rect 6097 1972 6099 1978
rect 6061 1944 6099 1972
rect 6133 1972 6135 1978
rect 6169 1978 6206 2006
rect 6169 1972 6171 1978
rect 6133 1944 6171 1972
rect 6205 1944 6206 1978
rect 6026 1938 6206 1944
rect 6026 1904 6063 1938
rect 6097 1904 6135 1938
rect 6169 1904 6206 1938
rect 6026 1870 6027 1904
rect 6061 1870 6099 1904
rect 6133 1870 6171 1904
rect 6205 1870 6206 1904
rect 6026 1836 6063 1870
rect 6097 1836 6135 1870
rect 6169 1836 6206 1870
rect 6026 1830 6206 1836
rect 6026 1796 6027 1830
rect 6061 1802 6099 1830
rect 6061 1796 6063 1802
rect 6026 1768 6063 1796
rect 6097 1796 6099 1802
rect 6133 1802 6171 1830
rect 6133 1796 6135 1802
rect 6097 1768 6135 1796
rect 6169 1796 6171 1802
rect 6205 1796 6206 1830
rect 6169 1768 6206 1796
rect 6026 1756 6206 1768
rect 6026 1722 6027 1756
rect 6061 1734 6099 1756
rect 6061 1722 6063 1734
rect 6026 1700 6063 1722
rect 6097 1722 6099 1734
rect 6133 1734 6171 1756
rect 6133 1722 6135 1734
rect 6097 1700 6135 1722
rect 6169 1722 6171 1734
rect 6205 1722 6206 1756
rect 6169 1700 6206 1722
rect 6026 1682 6206 1700
rect 6026 1648 6027 1682
rect 6061 1666 6099 1682
rect 6061 1648 6063 1666
rect 6026 1632 6063 1648
rect 6097 1648 6099 1666
rect 6133 1666 6171 1682
rect 6133 1648 6135 1666
rect 6097 1632 6135 1648
rect 6169 1648 6171 1666
rect 6205 1648 6206 1682
rect 6169 1632 6206 1648
rect 6026 1608 6206 1632
rect 6026 1574 6027 1608
rect 6061 1598 6099 1608
rect 6061 1574 6063 1598
rect 6026 1564 6063 1574
rect 6097 1574 6099 1598
rect 6133 1598 6171 1608
rect 6133 1574 6135 1598
rect 6097 1564 6135 1574
rect 6169 1574 6171 1598
rect 6205 1574 6206 1608
rect 6169 1564 6206 1574
rect 6026 1548 6206 1564
rect 6271 3104 6391 4200
rect 6833 4308 6953 4324
rect 6833 4274 6876 4308
rect 6910 4274 6953 4308
rect 6833 4234 6953 4274
rect 6833 4200 6876 4234
rect 6910 4200 6953 4234
rect 6271 3070 6314 3104
rect 6348 3070 6391 3104
rect 6271 3026 6391 3070
rect 6271 2992 6314 3026
rect 6348 2992 6391 3026
rect 6271 2948 6391 2992
rect 6271 2914 6314 2948
rect 6348 2914 6391 2948
rect 6271 2870 6391 2914
rect 6271 2836 6314 2870
rect 6348 2836 6391 2870
rect 6271 2792 6391 2836
rect 6271 2758 6314 2792
rect 6348 2758 6391 2792
rect 6271 2713 6391 2758
rect 6271 2679 6314 2713
rect 6348 2679 6391 2713
rect 6271 2634 6391 2679
rect 6271 2600 6314 2634
rect 6348 2600 6391 2634
rect 5841 1470 5884 1504
rect 5918 1470 5961 1504
rect 5841 1430 5961 1470
rect 5841 1396 5884 1430
rect 5918 1396 5961 1430
rect 5841 1250 5961 1396
rect 5841 1144 5848 1250
rect 5954 1144 5961 1250
rect 6271 1504 6391 2600
rect 6493 4092 6595 4118
rect 6629 4092 6731 4118
rect 6493 4082 6523 4092
rect 6701 4082 6731 4092
rect 6493 4014 6523 4048
rect 6701 4014 6731 4048
rect 6493 3946 6523 3980
rect 6701 3946 6731 3980
rect 6493 3878 6523 3912
rect 6701 3878 6731 3912
rect 6493 3810 6523 3844
rect 6701 3810 6731 3844
rect 6493 3742 6523 3776
rect 6701 3742 6731 3776
rect 6493 3674 6523 3708
rect 6701 3674 6731 3708
rect 6493 3606 6523 3640
rect 6701 3606 6731 3640
rect 6493 3538 6523 3572
rect 6701 3538 6731 3572
rect 6493 3470 6523 3504
rect 6701 3470 6731 3504
rect 6493 3402 6523 3436
rect 6701 3402 6731 3436
rect 6493 3334 6523 3368
rect 6701 3334 6731 3368
rect 6493 3266 6523 3300
rect 6701 3266 6731 3300
rect 6493 3198 6523 3232
rect 6701 3198 6731 3232
rect 6527 3164 6595 3194
rect 6629 3164 6697 3194
rect 6493 3148 6595 3164
rect 6629 3148 6731 3164
rect 6493 3108 6731 3148
rect 6493 3074 6523 3108
rect 6557 3074 6595 3108
rect 6629 3074 6667 3108
rect 6701 3074 6731 3108
rect 6493 3044 6731 3074
rect 6493 3028 6561 3044
rect 6493 2994 6523 3028
rect 6557 3010 6561 3028
rect 6595 3028 6629 3044
rect 6557 2994 6595 3010
rect 6663 3028 6731 3044
rect 6663 3010 6667 3028
rect 6629 2994 6667 3010
rect 6701 2994 6731 3028
rect 6493 2974 6731 2994
rect 6493 2948 6561 2974
rect 6493 2914 6523 2948
rect 6557 2940 6561 2948
rect 6595 2948 6629 2974
rect 6557 2914 6595 2940
rect 6663 2948 6731 2974
rect 6663 2940 6667 2948
rect 6629 2914 6667 2940
rect 6701 2914 6731 2948
rect 6493 2904 6731 2914
rect 6493 2870 6561 2904
rect 6595 2870 6629 2904
rect 6663 2870 6731 2904
rect 6493 2868 6731 2870
rect 6493 2834 6523 2868
rect 6557 2834 6595 2868
rect 6629 2834 6667 2868
rect 6701 2834 6731 2868
rect 6493 2800 6561 2834
rect 6595 2800 6629 2834
rect 6663 2800 6731 2834
rect 6493 2788 6731 2800
rect 6493 2754 6523 2788
rect 6557 2764 6595 2788
rect 6557 2754 6561 2764
rect 6493 2730 6561 2754
rect 6629 2764 6667 2788
rect 6595 2730 6629 2754
rect 6663 2754 6667 2764
rect 6701 2754 6731 2788
rect 6663 2730 6731 2754
rect 6493 2708 6731 2730
rect 6493 2674 6523 2708
rect 6557 2694 6595 2708
rect 6557 2674 6561 2694
rect 6493 2660 6561 2674
rect 6629 2694 6667 2708
rect 6595 2660 6629 2674
rect 6663 2674 6667 2694
rect 6701 2674 6731 2708
rect 6663 2660 6731 2674
rect 6493 2628 6731 2660
rect 6493 2594 6523 2628
rect 6557 2594 6595 2628
rect 6629 2594 6667 2628
rect 6701 2594 6731 2628
rect 6493 2556 6731 2594
rect 6493 2540 6595 2556
rect 6629 2540 6731 2556
rect 6527 2518 6595 2540
rect 6629 2518 6697 2540
rect 6493 2472 6523 2506
rect 6701 2472 6731 2506
rect 6493 2404 6523 2438
rect 6701 2404 6731 2438
rect 6493 2336 6523 2370
rect 6701 2336 6731 2370
rect 6493 2268 6523 2302
rect 6701 2268 6731 2302
rect 6493 2200 6523 2234
rect 6701 2200 6731 2234
rect 6493 2132 6523 2166
rect 6701 2132 6731 2166
rect 6493 2064 6523 2098
rect 6701 2064 6731 2098
rect 6493 1996 6523 2030
rect 6701 1996 6731 2030
rect 6493 1928 6523 1962
rect 6701 1928 6731 1962
rect 6493 1860 6523 1894
rect 6701 1860 6731 1894
rect 6493 1792 6523 1826
rect 6701 1792 6731 1826
rect 6493 1724 6523 1758
rect 6701 1724 6731 1758
rect 6493 1656 6523 1690
rect 6701 1656 6731 1690
rect 6493 1620 6523 1622
rect 6701 1620 6731 1622
rect 6493 1586 6595 1620
rect 6629 1586 6731 1620
rect 6493 1536 6731 1586
rect 6833 3104 6953 4200
rect 7263 4308 7383 4324
rect 7263 4274 7306 4308
rect 7340 4274 7383 4308
rect 7263 4234 7383 4274
rect 7263 4200 7306 4234
rect 7340 4200 7383 4234
rect 6833 3070 6876 3104
rect 6910 3070 6953 3104
rect 6833 3026 6953 3070
rect 6833 2992 6876 3026
rect 6910 2992 6953 3026
rect 6833 2948 6953 2992
rect 6833 2914 6876 2948
rect 6910 2914 6953 2948
rect 6833 2870 6953 2914
rect 6833 2836 6876 2870
rect 6910 2836 6953 2870
rect 6833 2792 6953 2836
rect 6833 2758 6876 2792
rect 6910 2758 6953 2792
rect 6833 2713 6953 2758
rect 6833 2679 6876 2713
rect 6910 2679 6953 2713
rect 6833 2634 6953 2679
rect 6833 2600 6876 2634
rect 6910 2600 6953 2634
rect 6271 1470 6314 1504
rect 6348 1470 6391 1504
rect 6271 1430 6391 1470
rect 6271 1396 6314 1430
rect 6348 1396 6391 1430
rect 6271 1250 6391 1396
rect 6271 1144 6278 1250
rect 6384 1144 6391 1250
rect 6833 1504 6953 2600
rect 7018 4064 7019 4098
rect 7053 4082 7091 4098
rect 7053 4064 7055 4082
rect 7018 4048 7055 4064
rect 7089 4064 7091 4082
rect 7125 4082 7163 4098
rect 7125 4064 7127 4082
rect 7089 4048 7127 4064
rect 7161 4064 7163 4082
rect 7197 4064 7198 4098
rect 7161 4048 7198 4064
rect 7018 4025 7198 4048
rect 7018 3991 7019 4025
rect 7053 4014 7091 4025
rect 7053 3991 7055 4014
rect 7018 3980 7055 3991
rect 7089 3991 7091 4014
rect 7125 4014 7163 4025
rect 7125 3991 7127 4014
rect 7089 3980 7127 3991
rect 7161 3991 7163 4014
rect 7197 3991 7198 4025
rect 7161 3980 7198 3991
rect 7018 3952 7198 3980
rect 7018 3918 7019 3952
rect 7053 3946 7091 3952
rect 7053 3918 7055 3946
rect 7018 3912 7055 3918
rect 7089 3918 7091 3946
rect 7125 3946 7163 3952
rect 7125 3918 7127 3946
rect 7089 3912 7127 3918
rect 7161 3918 7163 3946
rect 7197 3918 7198 3952
rect 7161 3912 7198 3918
rect 7018 3879 7198 3912
rect 7018 3845 7019 3879
rect 7053 3878 7091 3879
rect 7053 3845 7055 3878
rect 7018 3844 7055 3845
rect 7089 3845 7091 3878
rect 7125 3878 7163 3879
rect 7125 3845 7127 3878
rect 7089 3844 7127 3845
rect 7161 3845 7163 3878
rect 7197 3845 7198 3879
rect 7161 3844 7198 3845
rect 7018 3810 7198 3844
rect 7018 3806 7055 3810
rect 7018 3772 7019 3806
rect 7053 3776 7055 3806
rect 7089 3806 7127 3810
rect 7089 3776 7091 3806
rect 7053 3772 7091 3776
rect 7125 3776 7127 3806
rect 7161 3806 7198 3810
rect 7161 3776 7163 3806
rect 7125 3772 7163 3776
rect 7197 3772 7198 3806
rect 7018 3742 7198 3772
rect 7018 3733 7055 3742
rect 7018 3699 7019 3733
rect 7053 3708 7055 3733
rect 7089 3733 7127 3742
rect 7089 3708 7091 3733
rect 7053 3699 7091 3708
rect 7125 3708 7127 3733
rect 7161 3733 7198 3742
rect 7161 3708 7163 3733
rect 7125 3699 7163 3708
rect 7197 3699 7198 3733
rect 7018 3674 7198 3699
rect 7018 3660 7055 3674
rect 7018 3626 7019 3660
rect 7053 3640 7055 3660
rect 7089 3660 7127 3674
rect 7089 3640 7091 3660
rect 7053 3626 7091 3640
rect 7125 3640 7127 3660
rect 7161 3660 7198 3674
rect 7161 3640 7163 3660
rect 7125 3626 7163 3640
rect 7197 3626 7198 3660
rect 7018 3606 7198 3626
rect 7018 3587 7055 3606
rect 7018 3553 7019 3587
rect 7053 3572 7055 3587
rect 7089 3587 7127 3606
rect 7089 3572 7091 3587
rect 7053 3553 7091 3572
rect 7125 3572 7127 3587
rect 7161 3587 7198 3606
rect 7161 3572 7163 3587
rect 7125 3553 7163 3572
rect 7197 3553 7198 3587
rect 7018 3538 7198 3553
rect 7018 3514 7055 3538
rect 7018 3480 7019 3514
rect 7053 3504 7055 3514
rect 7089 3514 7127 3538
rect 7089 3504 7091 3514
rect 7053 3480 7091 3504
rect 7125 3504 7127 3514
rect 7161 3514 7198 3538
rect 7161 3504 7163 3514
rect 7125 3480 7163 3504
rect 7197 3480 7198 3514
rect 7018 3470 7198 3480
rect 7018 3441 7055 3470
rect 7018 3407 7019 3441
rect 7053 3436 7055 3441
rect 7089 3441 7127 3470
rect 7089 3436 7091 3441
rect 7053 3407 7091 3436
rect 7125 3436 7127 3441
rect 7161 3441 7198 3470
rect 7161 3436 7163 3441
rect 7125 3407 7163 3436
rect 7197 3407 7198 3441
rect 7018 3402 7198 3407
rect 7018 3368 7055 3402
rect 7089 3368 7127 3402
rect 7161 3368 7198 3402
rect 7018 3334 7019 3368
rect 7053 3334 7091 3368
rect 7125 3334 7163 3368
rect 7197 3334 7198 3368
rect 7018 3300 7055 3334
rect 7089 3300 7127 3334
rect 7161 3300 7198 3334
rect 7018 3295 7198 3300
rect 7018 3261 7019 3295
rect 7053 3266 7091 3295
rect 7053 3261 7055 3266
rect 7018 3232 7055 3261
rect 7089 3261 7091 3266
rect 7125 3266 7163 3295
rect 7125 3261 7127 3266
rect 7089 3232 7127 3261
rect 7161 3261 7163 3266
rect 7197 3261 7198 3295
rect 7161 3232 7198 3261
rect 7018 3222 7198 3232
rect 7018 3188 7019 3222
rect 7053 3198 7091 3222
rect 7053 3188 7055 3198
rect 7018 3164 7055 3188
rect 7089 3188 7091 3198
rect 7125 3198 7163 3222
rect 7125 3188 7127 3198
rect 7089 3164 7127 3188
rect 7161 3188 7163 3198
rect 7197 3188 7198 3222
rect 7161 3164 7198 3188
rect 7018 3149 7198 3164
rect 7018 3115 7019 3149
rect 7053 3115 7091 3149
rect 7125 3115 7163 3149
rect 7197 3115 7198 3149
rect 7018 3076 7198 3115
rect 7018 3042 7019 3076
rect 7053 3042 7091 3076
rect 7125 3042 7163 3076
rect 7197 3042 7198 3076
rect 7018 3003 7198 3042
rect 7018 2969 7019 3003
rect 7053 2969 7091 3003
rect 7125 2969 7163 3003
rect 7197 2969 7198 3003
rect 7018 2930 7198 2969
rect 7018 2896 7019 2930
rect 7053 2896 7091 2930
rect 7125 2896 7163 2930
rect 7197 2896 7198 2930
rect 7018 2857 7198 2896
rect 7018 2823 7019 2857
rect 7053 2823 7091 2857
rect 7125 2823 7163 2857
rect 7197 2823 7198 2857
rect 7018 2784 7198 2823
rect 7018 2750 7019 2784
rect 7053 2750 7091 2784
rect 7125 2750 7163 2784
rect 7197 2750 7198 2784
rect 7018 2711 7198 2750
rect 7018 2677 7019 2711
rect 7053 2677 7091 2711
rect 7125 2677 7163 2711
rect 7197 2677 7198 2711
rect 7018 2638 7198 2677
rect 7018 2604 7019 2638
rect 7053 2604 7091 2638
rect 7125 2604 7163 2638
rect 7197 2604 7198 2638
rect 7018 2565 7198 2604
rect 7018 2531 7019 2565
rect 7053 2531 7091 2565
rect 7125 2531 7163 2565
rect 7197 2531 7198 2565
rect 7018 2492 7198 2531
rect 7018 2458 7019 2492
rect 7053 2482 7091 2492
rect 7053 2458 7055 2482
rect 7018 2448 7055 2458
rect 7089 2458 7091 2482
rect 7125 2482 7163 2492
rect 7125 2458 7127 2482
rect 7089 2448 7127 2458
rect 7161 2458 7163 2482
rect 7197 2458 7198 2492
rect 7161 2448 7198 2458
rect 7018 2419 7198 2448
rect 7018 2385 7019 2419
rect 7053 2414 7091 2419
rect 7053 2385 7055 2414
rect 7018 2380 7055 2385
rect 7089 2385 7091 2414
rect 7125 2414 7163 2419
rect 7125 2385 7127 2414
rect 7089 2380 7127 2385
rect 7161 2385 7163 2414
rect 7197 2385 7198 2419
rect 7161 2380 7198 2385
rect 7018 2346 7198 2380
rect 7018 2312 7019 2346
rect 7053 2312 7055 2346
rect 7089 2312 7091 2346
rect 7125 2312 7127 2346
rect 7161 2312 7163 2346
rect 7197 2312 7198 2346
rect 7018 2278 7198 2312
rect 7018 2273 7055 2278
rect 7018 2239 7019 2273
rect 7053 2244 7055 2273
rect 7089 2273 7127 2278
rect 7089 2244 7091 2273
rect 7053 2239 7091 2244
rect 7125 2244 7127 2273
rect 7161 2273 7198 2278
rect 7161 2244 7163 2273
rect 7125 2239 7163 2244
rect 7197 2239 7198 2273
rect 7018 2210 7198 2239
rect 7018 2200 7055 2210
rect 7018 2166 7019 2200
rect 7053 2176 7055 2200
rect 7089 2200 7127 2210
rect 7089 2176 7091 2200
rect 7053 2166 7091 2176
rect 7125 2176 7127 2200
rect 7161 2200 7198 2210
rect 7161 2176 7163 2200
rect 7125 2166 7163 2176
rect 7197 2166 7198 2200
rect 7018 2142 7198 2166
rect 7018 2126 7055 2142
rect 7018 2092 7019 2126
rect 7053 2108 7055 2126
rect 7089 2126 7127 2142
rect 7089 2108 7091 2126
rect 7053 2092 7091 2108
rect 7125 2108 7127 2126
rect 7161 2126 7198 2142
rect 7161 2108 7163 2126
rect 7125 2092 7163 2108
rect 7197 2092 7198 2126
rect 7018 2074 7198 2092
rect 7018 2052 7055 2074
rect 7018 2018 7019 2052
rect 7053 2040 7055 2052
rect 7089 2052 7127 2074
rect 7089 2040 7091 2052
rect 7053 2018 7091 2040
rect 7125 2040 7127 2052
rect 7161 2052 7198 2074
rect 7161 2040 7163 2052
rect 7125 2018 7163 2040
rect 7197 2018 7198 2052
rect 7018 2006 7198 2018
rect 7018 1978 7055 2006
rect 7018 1944 7019 1978
rect 7053 1972 7055 1978
rect 7089 1978 7127 2006
rect 7089 1972 7091 1978
rect 7053 1944 7091 1972
rect 7125 1972 7127 1978
rect 7161 1978 7198 2006
rect 7161 1972 7163 1978
rect 7125 1944 7163 1972
rect 7197 1944 7198 1978
rect 7018 1938 7198 1944
rect 7018 1904 7055 1938
rect 7089 1904 7127 1938
rect 7161 1904 7198 1938
rect 7018 1870 7019 1904
rect 7053 1870 7091 1904
rect 7125 1870 7163 1904
rect 7197 1870 7198 1904
rect 7018 1836 7055 1870
rect 7089 1836 7127 1870
rect 7161 1836 7198 1870
rect 7018 1830 7198 1836
rect 7018 1796 7019 1830
rect 7053 1802 7091 1830
rect 7053 1796 7055 1802
rect 7018 1768 7055 1796
rect 7089 1796 7091 1802
rect 7125 1802 7163 1830
rect 7125 1796 7127 1802
rect 7089 1768 7127 1796
rect 7161 1796 7163 1802
rect 7197 1796 7198 1830
rect 7161 1768 7198 1796
rect 7018 1756 7198 1768
rect 7018 1722 7019 1756
rect 7053 1734 7091 1756
rect 7053 1722 7055 1734
rect 7018 1700 7055 1722
rect 7089 1722 7091 1734
rect 7125 1734 7163 1756
rect 7125 1722 7127 1734
rect 7089 1700 7127 1722
rect 7161 1722 7163 1734
rect 7197 1722 7198 1756
rect 7161 1700 7198 1722
rect 7018 1682 7198 1700
rect 7018 1648 7019 1682
rect 7053 1666 7091 1682
rect 7053 1648 7055 1666
rect 7018 1632 7055 1648
rect 7089 1648 7091 1666
rect 7125 1666 7163 1682
rect 7125 1648 7127 1666
rect 7089 1632 7127 1648
rect 7161 1648 7163 1666
rect 7197 1648 7198 1682
rect 7161 1632 7198 1648
rect 7018 1608 7198 1632
rect 7018 1574 7019 1608
rect 7053 1598 7091 1608
rect 7053 1574 7055 1598
rect 7018 1564 7055 1574
rect 7089 1574 7091 1598
rect 7125 1598 7163 1608
rect 7125 1574 7127 1598
rect 7089 1564 7127 1574
rect 7161 1574 7163 1598
rect 7197 1574 7198 1608
rect 7161 1564 7198 1574
rect 7018 1548 7198 1564
rect 7263 3104 7383 4200
rect 7825 4308 7945 4324
rect 7825 4274 7868 4308
rect 7902 4274 7945 4308
rect 7825 4234 7945 4274
rect 7825 4200 7868 4234
rect 7902 4200 7945 4234
rect 7263 3070 7306 3104
rect 7340 3070 7383 3104
rect 7263 3026 7383 3070
rect 7263 2992 7306 3026
rect 7340 2992 7383 3026
rect 7263 2948 7383 2992
rect 7263 2914 7306 2948
rect 7340 2914 7383 2948
rect 7263 2870 7383 2914
rect 7263 2836 7306 2870
rect 7340 2836 7383 2870
rect 7263 2792 7383 2836
rect 7263 2758 7306 2792
rect 7340 2758 7383 2792
rect 7263 2713 7383 2758
rect 7263 2679 7306 2713
rect 7340 2679 7383 2713
rect 7263 2634 7383 2679
rect 7263 2600 7306 2634
rect 7340 2600 7383 2634
rect 6833 1470 6876 1504
rect 6910 1470 6953 1504
rect 6833 1430 6953 1470
rect 6833 1396 6876 1430
rect 6910 1396 6953 1430
rect 6833 1250 6953 1396
rect 6833 1144 6840 1250
rect 6946 1144 6953 1250
rect 7263 1504 7383 2600
rect 7485 4092 7587 4118
rect 7621 4092 7723 4118
rect 7485 4082 7515 4092
rect 7693 4082 7723 4092
rect 7485 4014 7515 4048
rect 7693 4014 7723 4048
rect 7485 3946 7515 3980
rect 7693 3946 7723 3980
rect 7485 3878 7515 3912
rect 7693 3878 7723 3912
rect 7485 3810 7515 3844
rect 7693 3810 7723 3844
rect 7485 3742 7515 3776
rect 7693 3742 7723 3776
rect 7485 3674 7515 3708
rect 7693 3674 7723 3708
rect 7485 3606 7515 3640
rect 7693 3606 7723 3640
rect 7485 3538 7515 3572
rect 7693 3538 7723 3572
rect 7485 3470 7515 3504
rect 7693 3470 7723 3504
rect 7485 3402 7515 3436
rect 7693 3402 7723 3436
rect 7485 3334 7515 3368
rect 7693 3334 7723 3368
rect 7485 3266 7515 3300
rect 7693 3266 7723 3300
rect 7485 3198 7515 3232
rect 7693 3198 7723 3232
rect 7519 3164 7587 3194
rect 7621 3164 7689 3194
rect 7485 3148 7587 3164
rect 7621 3148 7723 3164
rect 7485 3108 7723 3148
rect 7485 3074 7515 3108
rect 7549 3074 7587 3108
rect 7621 3074 7659 3108
rect 7693 3074 7723 3108
rect 7485 3044 7723 3074
rect 7485 3028 7553 3044
rect 7485 2994 7515 3028
rect 7549 3010 7553 3028
rect 7587 3028 7621 3044
rect 7549 2994 7587 3010
rect 7655 3028 7723 3044
rect 7655 3010 7659 3028
rect 7621 2994 7659 3010
rect 7693 2994 7723 3028
rect 7485 2974 7723 2994
rect 7485 2948 7553 2974
rect 7485 2914 7515 2948
rect 7549 2940 7553 2948
rect 7587 2948 7621 2974
rect 7549 2914 7587 2940
rect 7655 2948 7723 2974
rect 7655 2940 7659 2948
rect 7621 2914 7659 2940
rect 7693 2914 7723 2948
rect 7485 2904 7723 2914
rect 7485 2870 7553 2904
rect 7587 2870 7621 2904
rect 7655 2870 7723 2904
rect 7485 2868 7723 2870
rect 7485 2834 7515 2868
rect 7549 2834 7587 2868
rect 7621 2834 7659 2868
rect 7693 2834 7723 2868
rect 7485 2800 7553 2834
rect 7587 2800 7621 2834
rect 7655 2800 7723 2834
rect 7485 2788 7723 2800
rect 7485 2754 7515 2788
rect 7549 2764 7587 2788
rect 7549 2754 7553 2764
rect 7485 2730 7553 2754
rect 7621 2764 7659 2788
rect 7587 2730 7621 2754
rect 7655 2754 7659 2764
rect 7693 2754 7723 2788
rect 7655 2730 7723 2754
rect 7485 2708 7723 2730
rect 7485 2674 7515 2708
rect 7549 2694 7587 2708
rect 7549 2674 7553 2694
rect 7485 2660 7553 2674
rect 7621 2694 7659 2708
rect 7587 2660 7621 2674
rect 7655 2674 7659 2694
rect 7693 2674 7723 2708
rect 7655 2660 7723 2674
rect 7485 2628 7723 2660
rect 7485 2594 7515 2628
rect 7549 2594 7587 2628
rect 7621 2594 7659 2628
rect 7693 2594 7723 2628
rect 7485 2556 7723 2594
rect 7485 2540 7587 2556
rect 7621 2540 7723 2556
rect 7519 2518 7587 2540
rect 7621 2518 7689 2540
rect 7485 2472 7515 2506
rect 7693 2472 7723 2506
rect 7485 2404 7515 2438
rect 7693 2404 7723 2438
rect 7485 2336 7515 2370
rect 7693 2336 7723 2370
rect 7485 2268 7515 2302
rect 7693 2268 7723 2302
rect 7485 2200 7515 2234
rect 7693 2200 7723 2234
rect 7485 2132 7515 2166
rect 7693 2132 7723 2166
rect 7485 2064 7515 2098
rect 7693 2064 7723 2098
rect 7485 1996 7515 2030
rect 7693 1996 7723 2030
rect 7485 1928 7515 1962
rect 7693 1928 7723 1962
rect 7485 1860 7515 1894
rect 7693 1860 7723 1894
rect 7485 1792 7515 1826
rect 7693 1792 7723 1826
rect 7485 1724 7515 1758
rect 7693 1724 7723 1758
rect 7485 1656 7515 1690
rect 7693 1656 7723 1690
rect 7485 1620 7515 1622
rect 7693 1620 7723 1622
rect 7485 1586 7587 1620
rect 7621 1586 7723 1620
rect 7485 1536 7723 1586
rect 7825 3104 7945 4200
rect 8255 4308 8375 4324
rect 8255 4274 8298 4308
rect 8332 4274 8375 4308
rect 8255 4234 8375 4274
rect 8255 4200 8298 4234
rect 8332 4200 8375 4234
rect 7825 3070 7868 3104
rect 7902 3070 7945 3104
rect 7825 3026 7945 3070
rect 7825 2992 7868 3026
rect 7902 2992 7945 3026
rect 7825 2948 7945 2992
rect 7825 2914 7868 2948
rect 7902 2914 7945 2948
rect 7825 2870 7945 2914
rect 7825 2836 7868 2870
rect 7902 2836 7945 2870
rect 7825 2792 7945 2836
rect 7825 2758 7868 2792
rect 7902 2758 7945 2792
rect 7825 2713 7945 2758
rect 7825 2679 7868 2713
rect 7902 2679 7945 2713
rect 7825 2634 7945 2679
rect 7825 2600 7868 2634
rect 7902 2600 7945 2634
rect 7263 1470 7306 1504
rect 7340 1470 7383 1504
rect 7263 1430 7383 1470
rect 7263 1396 7306 1430
rect 7340 1396 7383 1430
rect 7263 1250 7383 1396
rect 7263 1144 7270 1250
rect 7376 1144 7383 1250
rect 7825 1504 7945 2600
rect 8010 4064 8011 4098
rect 8045 4082 8083 4098
rect 8045 4064 8047 4082
rect 8010 4048 8047 4064
rect 8081 4064 8083 4082
rect 8117 4082 8155 4098
rect 8117 4064 8119 4082
rect 8081 4048 8119 4064
rect 8153 4064 8155 4082
rect 8189 4064 8190 4098
rect 8153 4048 8190 4064
rect 8010 4025 8190 4048
rect 8010 3991 8011 4025
rect 8045 4014 8083 4025
rect 8045 3991 8047 4014
rect 8010 3980 8047 3991
rect 8081 3991 8083 4014
rect 8117 4014 8155 4025
rect 8117 3991 8119 4014
rect 8081 3980 8119 3991
rect 8153 3991 8155 4014
rect 8189 3991 8190 4025
rect 8153 3980 8190 3991
rect 8010 3952 8190 3980
rect 8010 3918 8011 3952
rect 8045 3946 8083 3952
rect 8045 3918 8047 3946
rect 8010 3912 8047 3918
rect 8081 3918 8083 3946
rect 8117 3946 8155 3952
rect 8117 3918 8119 3946
rect 8081 3912 8119 3918
rect 8153 3918 8155 3946
rect 8189 3918 8190 3952
rect 8153 3912 8190 3918
rect 8010 3879 8190 3912
rect 8010 3845 8011 3879
rect 8045 3878 8083 3879
rect 8045 3845 8047 3878
rect 8010 3844 8047 3845
rect 8081 3845 8083 3878
rect 8117 3878 8155 3879
rect 8117 3845 8119 3878
rect 8081 3844 8119 3845
rect 8153 3845 8155 3878
rect 8189 3845 8190 3879
rect 8153 3844 8190 3845
rect 8010 3810 8190 3844
rect 8010 3806 8047 3810
rect 8010 3772 8011 3806
rect 8045 3776 8047 3806
rect 8081 3806 8119 3810
rect 8081 3776 8083 3806
rect 8045 3772 8083 3776
rect 8117 3776 8119 3806
rect 8153 3806 8190 3810
rect 8153 3776 8155 3806
rect 8117 3772 8155 3776
rect 8189 3772 8190 3806
rect 8010 3742 8190 3772
rect 8010 3733 8047 3742
rect 8010 3699 8011 3733
rect 8045 3708 8047 3733
rect 8081 3733 8119 3742
rect 8081 3708 8083 3733
rect 8045 3699 8083 3708
rect 8117 3708 8119 3733
rect 8153 3733 8190 3742
rect 8153 3708 8155 3733
rect 8117 3699 8155 3708
rect 8189 3699 8190 3733
rect 8010 3674 8190 3699
rect 8010 3660 8047 3674
rect 8010 3626 8011 3660
rect 8045 3640 8047 3660
rect 8081 3660 8119 3674
rect 8081 3640 8083 3660
rect 8045 3626 8083 3640
rect 8117 3640 8119 3660
rect 8153 3660 8190 3674
rect 8153 3640 8155 3660
rect 8117 3626 8155 3640
rect 8189 3626 8190 3660
rect 8010 3606 8190 3626
rect 8010 3587 8047 3606
rect 8010 3553 8011 3587
rect 8045 3572 8047 3587
rect 8081 3587 8119 3606
rect 8081 3572 8083 3587
rect 8045 3553 8083 3572
rect 8117 3572 8119 3587
rect 8153 3587 8190 3606
rect 8153 3572 8155 3587
rect 8117 3553 8155 3572
rect 8189 3553 8190 3587
rect 8010 3538 8190 3553
rect 8010 3514 8047 3538
rect 8010 3480 8011 3514
rect 8045 3504 8047 3514
rect 8081 3514 8119 3538
rect 8081 3504 8083 3514
rect 8045 3480 8083 3504
rect 8117 3504 8119 3514
rect 8153 3514 8190 3538
rect 8153 3504 8155 3514
rect 8117 3480 8155 3504
rect 8189 3480 8190 3514
rect 8010 3470 8190 3480
rect 8010 3441 8047 3470
rect 8010 3407 8011 3441
rect 8045 3436 8047 3441
rect 8081 3441 8119 3470
rect 8081 3436 8083 3441
rect 8045 3407 8083 3436
rect 8117 3436 8119 3441
rect 8153 3441 8190 3470
rect 8153 3436 8155 3441
rect 8117 3407 8155 3436
rect 8189 3407 8190 3441
rect 8010 3402 8190 3407
rect 8010 3368 8047 3402
rect 8081 3368 8119 3402
rect 8153 3368 8190 3402
rect 8010 3334 8011 3368
rect 8045 3334 8083 3368
rect 8117 3334 8155 3368
rect 8189 3334 8190 3368
rect 8010 3300 8047 3334
rect 8081 3300 8119 3334
rect 8153 3300 8190 3334
rect 8010 3295 8190 3300
rect 8010 3261 8011 3295
rect 8045 3266 8083 3295
rect 8045 3261 8047 3266
rect 8010 3232 8047 3261
rect 8081 3261 8083 3266
rect 8117 3266 8155 3295
rect 8117 3261 8119 3266
rect 8081 3232 8119 3261
rect 8153 3261 8155 3266
rect 8189 3261 8190 3295
rect 8153 3232 8190 3261
rect 8010 3222 8190 3232
rect 8010 3188 8011 3222
rect 8045 3198 8083 3222
rect 8045 3188 8047 3198
rect 8010 3164 8047 3188
rect 8081 3188 8083 3198
rect 8117 3198 8155 3222
rect 8117 3188 8119 3198
rect 8081 3164 8119 3188
rect 8153 3188 8155 3198
rect 8189 3188 8190 3222
rect 8153 3164 8190 3188
rect 8010 3149 8190 3164
rect 8010 3115 8011 3149
rect 8045 3115 8083 3149
rect 8117 3115 8155 3149
rect 8189 3115 8190 3149
rect 8010 3076 8190 3115
rect 8010 3042 8011 3076
rect 8045 3042 8083 3076
rect 8117 3042 8155 3076
rect 8189 3042 8190 3076
rect 8010 3003 8190 3042
rect 8010 2969 8011 3003
rect 8045 2969 8083 3003
rect 8117 2969 8155 3003
rect 8189 2969 8190 3003
rect 8010 2930 8190 2969
rect 8010 2896 8011 2930
rect 8045 2896 8083 2930
rect 8117 2896 8155 2930
rect 8189 2896 8190 2930
rect 8010 2857 8190 2896
rect 8010 2823 8011 2857
rect 8045 2823 8083 2857
rect 8117 2823 8155 2857
rect 8189 2823 8190 2857
rect 8010 2784 8190 2823
rect 8010 2750 8011 2784
rect 8045 2750 8083 2784
rect 8117 2750 8155 2784
rect 8189 2750 8190 2784
rect 8010 2711 8190 2750
rect 8010 2677 8011 2711
rect 8045 2677 8083 2711
rect 8117 2677 8155 2711
rect 8189 2677 8190 2711
rect 8010 2638 8190 2677
rect 8010 2604 8011 2638
rect 8045 2604 8083 2638
rect 8117 2604 8155 2638
rect 8189 2604 8190 2638
rect 8010 2565 8190 2604
rect 8010 2531 8011 2565
rect 8045 2531 8083 2565
rect 8117 2531 8155 2565
rect 8189 2531 8190 2565
rect 8010 2492 8190 2531
rect 8010 2458 8011 2492
rect 8045 2482 8083 2492
rect 8045 2458 8047 2482
rect 8010 2448 8047 2458
rect 8081 2458 8083 2482
rect 8117 2482 8155 2492
rect 8117 2458 8119 2482
rect 8081 2448 8119 2458
rect 8153 2458 8155 2482
rect 8189 2458 8190 2492
rect 8153 2448 8190 2458
rect 8010 2419 8190 2448
rect 8010 2385 8011 2419
rect 8045 2414 8083 2419
rect 8045 2385 8047 2414
rect 8010 2380 8047 2385
rect 8081 2385 8083 2414
rect 8117 2414 8155 2419
rect 8117 2385 8119 2414
rect 8081 2380 8119 2385
rect 8153 2385 8155 2414
rect 8189 2385 8190 2419
rect 8153 2380 8190 2385
rect 8010 2346 8190 2380
rect 8010 2312 8011 2346
rect 8045 2312 8047 2346
rect 8081 2312 8083 2346
rect 8117 2312 8119 2346
rect 8153 2312 8155 2346
rect 8189 2312 8190 2346
rect 8010 2278 8190 2312
rect 8010 2273 8047 2278
rect 8010 2239 8011 2273
rect 8045 2244 8047 2273
rect 8081 2273 8119 2278
rect 8081 2244 8083 2273
rect 8045 2239 8083 2244
rect 8117 2244 8119 2273
rect 8153 2273 8190 2278
rect 8153 2244 8155 2273
rect 8117 2239 8155 2244
rect 8189 2239 8190 2273
rect 8010 2210 8190 2239
rect 8010 2200 8047 2210
rect 8010 2166 8011 2200
rect 8045 2176 8047 2200
rect 8081 2200 8119 2210
rect 8081 2176 8083 2200
rect 8045 2166 8083 2176
rect 8117 2176 8119 2200
rect 8153 2200 8190 2210
rect 8153 2176 8155 2200
rect 8117 2166 8155 2176
rect 8189 2166 8190 2200
rect 8010 2142 8190 2166
rect 8010 2126 8047 2142
rect 8010 2092 8011 2126
rect 8045 2108 8047 2126
rect 8081 2126 8119 2142
rect 8081 2108 8083 2126
rect 8045 2092 8083 2108
rect 8117 2108 8119 2126
rect 8153 2126 8190 2142
rect 8153 2108 8155 2126
rect 8117 2092 8155 2108
rect 8189 2092 8190 2126
rect 8010 2074 8190 2092
rect 8010 2052 8047 2074
rect 8010 2018 8011 2052
rect 8045 2040 8047 2052
rect 8081 2052 8119 2074
rect 8081 2040 8083 2052
rect 8045 2018 8083 2040
rect 8117 2040 8119 2052
rect 8153 2052 8190 2074
rect 8153 2040 8155 2052
rect 8117 2018 8155 2040
rect 8189 2018 8190 2052
rect 8010 2006 8190 2018
rect 8010 1978 8047 2006
rect 8010 1944 8011 1978
rect 8045 1972 8047 1978
rect 8081 1978 8119 2006
rect 8081 1972 8083 1978
rect 8045 1944 8083 1972
rect 8117 1972 8119 1978
rect 8153 1978 8190 2006
rect 8153 1972 8155 1978
rect 8117 1944 8155 1972
rect 8189 1944 8190 1978
rect 8010 1938 8190 1944
rect 8010 1904 8047 1938
rect 8081 1904 8119 1938
rect 8153 1904 8190 1938
rect 8010 1870 8011 1904
rect 8045 1870 8083 1904
rect 8117 1870 8155 1904
rect 8189 1870 8190 1904
rect 8010 1836 8047 1870
rect 8081 1836 8119 1870
rect 8153 1836 8190 1870
rect 8010 1830 8190 1836
rect 8010 1796 8011 1830
rect 8045 1802 8083 1830
rect 8045 1796 8047 1802
rect 8010 1768 8047 1796
rect 8081 1796 8083 1802
rect 8117 1802 8155 1830
rect 8117 1796 8119 1802
rect 8081 1768 8119 1796
rect 8153 1796 8155 1802
rect 8189 1796 8190 1830
rect 8153 1768 8190 1796
rect 8010 1756 8190 1768
rect 8010 1722 8011 1756
rect 8045 1734 8083 1756
rect 8045 1722 8047 1734
rect 8010 1700 8047 1722
rect 8081 1722 8083 1734
rect 8117 1734 8155 1756
rect 8117 1722 8119 1734
rect 8081 1700 8119 1722
rect 8153 1722 8155 1734
rect 8189 1722 8190 1756
rect 8153 1700 8190 1722
rect 8010 1682 8190 1700
rect 8010 1648 8011 1682
rect 8045 1666 8083 1682
rect 8045 1648 8047 1666
rect 8010 1632 8047 1648
rect 8081 1648 8083 1666
rect 8117 1666 8155 1682
rect 8117 1648 8119 1666
rect 8081 1632 8119 1648
rect 8153 1648 8155 1666
rect 8189 1648 8190 1682
rect 8153 1632 8190 1648
rect 8010 1608 8190 1632
rect 8010 1574 8011 1608
rect 8045 1598 8083 1608
rect 8045 1574 8047 1598
rect 8010 1564 8047 1574
rect 8081 1574 8083 1598
rect 8117 1598 8155 1608
rect 8117 1574 8119 1598
rect 8081 1564 8119 1574
rect 8153 1574 8155 1598
rect 8189 1574 8190 1608
rect 8153 1564 8190 1574
rect 8010 1548 8190 1564
rect 8255 3104 8375 4200
rect 8817 4308 8937 4324
rect 8817 4274 8860 4308
rect 8894 4274 8937 4308
rect 8817 4234 8937 4274
rect 8817 4200 8860 4234
rect 8894 4200 8937 4234
rect 8255 3070 8298 3104
rect 8332 3070 8375 3104
rect 8255 3026 8375 3070
rect 8255 2992 8298 3026
rect 8332 2992 8375 3026
rect 8255 2948 8375 2992
rect 8255 2914 8298 2948
rect 8332 2914 8375 2948
rect 8255 2870 8375 2914
rect 8255 2836 8298 2870
rect 8332 2836 8375 2870
rect 8255 2792 8375 2836
rect 8255 2758 8298 2792
rect 8332 2758 8375 2792
rect 8255 2713 8375 2758
rect 8255 2679 8298 2713
rect 8332 2679 8375 2713
rect 8255 2634 8375 2679
rect 8255 2600 8298 2634
rect 8332 2600 8375 2634
rect 7825 1470 7868 1504
rect 7902 1470 7945 1504
rect 7825 1430 7945 1470
rect 7825 1396 7868 1430
rect 7902 1396 7945 1430
rect 7825 1250 7945 1396
rect 7825 1144 7832 1250
rect 7938 1144 7945 1250
rect 8255 1504 8375 2600
rect 8477 4092 8579 4118
rect 8613 4092 8715 4118
rect 8477 4082 8507 4092
rect 8685 4082 8715 4092
rect 8477 4014 8507 4048
rect 8685 4014 8715 4048
rect 8477 3946 8507 3980
rect 8685 3946 8715 3980
rect 8477 3878 8507 3912
rect 8685 3878 8715 3912
rect 8477 3810 8507 3844
rect 8685 3810 8715 3844
rect 8477 3742 8507 3776
rect 8685 3742 8715 3776
rect 8477 3674 8507 3708
rect 8685 3674 8715 3708
rect 8477 3606 8507 3640
rect 8685 3606 8715 3640
rect 8477 3538 8507 3572
rect 8685 3538 8715 3572
rect 8477 3470 8507 3504
rect 8685 3470 8715 3504
rect 8477 3402 8507 3436
rect 8685 3402 8715 3436
rect 8477 3334 8507 3368
rect 8685 3334 8715 3368
rect 8477 3266 8507 3300
rect 8685 3266 8715 3300
rect 8477 3198 8507 3232
rect 8685 3198 8715 3232
rect 8511 3164 8579 3194
rect 8613 3164 8681 3194
rect 8477 3148 8579 3164
rect 8613 3148 8715 3164
rect 8477 3108 8715 3148
rect 8477 3074 8507 3108
rect 8541 3074 8579 3108
rect 8613 3074 8651 3108
rect 8685 3074 8715 3108
rect 8477 3044 8715 3074
rect 8477 3028 8545 3044
rect 8477 2994 8507 3028
rect 8541 3010 8545 3028
rect 8579 3028 8613 3044
rect 8541 2994 8579 3010
rect 8647 3028 8715 3044
rect 8647 3010 8651 3028
rect 8613 2994 8651 3010
rect 8685 2994 8715 3028
rect 8477 2974 8715 2994
rect 8477 2948 8545 2974
rect 8477 2914 8507 2948
rect 8541 2940 8545 2948
rect 8579 2948 8613 2974
rect 8541 2914 8579 2940
rect 8647 2948 8715 2974
rect 8647 2940 8651 2948
rect 8613 2914 8651 2940
rect 8685 2914 8715 2948
rect 8477 2904 8715 2914
rect 8477 2870 8545 2904
rect 8579 2870 8613 2904
rect 8647 2870 8715 2904
rect 8477 2868 8715 2870
rect 8477 2834 8507 2868
rect 8541 2834 8579 2868
rect 8613 2834 8651 2868
rect 8685 2834 8715 2868
rect 8477 2800 8545 2834
rect 8579 2800 8613 2834
rect 8647 2800 8715 2834
rect 8477 2788 8715 2800
rect 8477 2754 8507 2788
rect 8541 2764 8579 2788
rect 8541 2754 8545 2764
rect 8477 2730 8545 2754
rect 8613 2764 8651 2788
rect 8579 2730 8613 2754
rect 8647 2754 8651 2764
rect 8685 2754 8715 2788
rect 8647 2730 8715 2754
rect 8477 2708 8715 2730
rect 8477 2674 8507 2708
rect 8541 2694 8579 2708
rect 8541 2674 8545 2694
rect 8477 2660 8545 2674
rect 8613 2694 8651 2708
rect 8579 2660 8613 2674
rect 8647 2674 8651 2694
rect 8685 2674 8715 2708
rect 8647 2660 8715 2674
rect 8477 2628 8715 2660
rect 8477 2594 8507 2628
rect 8541 2594 8579 2628
rect 8613 2594 8651 2628
rect 8685 2594 8715 2628
rect 8477 2556 8715 2594
rect 8477 2540 8579 2556
rect 8613 2540 8715 2556
rect 8511 2518 8579 2540
rect 8613 2518 8681 2540
rect 8477 2472 8507 2506
rect 8685 2472 8715 2506
rect 8477 2404 8507 2438
rect 8685 2404 8715 2438
rect 8477 2336 8507 2370
rect 8685 2336 8715 2370
rect 8477 2268 8507 2302
rect 8685 2268 8715 2302
rect 8477 2200 8507 2234
rect 8685 2200 8715 2234
rect 8477 2132 8507 2166
rect 8685 2132 8715 2166
rect 8477 2064 8507 2098
rect 8685 2064 8715 2098
rect 8477 1996 8507 2030
rect 8685 1996 8715 2030
rect 8477 1928 8507 1962
rect 8685 1928 8715 1962
rect 8477 1860 8507 1894
rect 8685 1860 8715 1894
rect 8477 1792 8507 1826
rect 8685 1792 8715 1826
rect 8477 1724 8507 1758
rect 8685 1724 8715 1758
rect 8477 1656 8507 1690
rect 8685 1656 8715 1690
rect 8477 1620 8507 1622
rect 8685 1620 8715 1622
rect 8477 1586 8579 1620
rect 8613 1586 8715 1620
rect 8477 1536 8715 1586
rect 8817 3104 8937 4200
rect 9247 4308 9367 4324
rect 9247 4274 9290 4308
rect 9324 4274 9367 4308
rect 9247 4234 9367 4274
rect 9247 4200 9290 4234
rect 9324 4200 9367 4234
rect 8817 3070 8860 3104
rect 8894 3070 8937 3104
rect 8817 3026 8937 3070
rect 8817 2992 8860 3026
rect 8894 2992 8937 3026
rect 8817 2948 8937 2992
rect 8817 2914 8860 2948
rect 8894 2914 8937 2948
rect 8817 2870 8937 2914
rect 8817 2836 8860 2870
rect 8894 2836 8937 2870
rect 8817 2792 8937 2836
rect 8817 2758 8860 2792
rect 8894 2758 8937 2792
rect 8817 2713 8937 2758
rect 8817 2679 8860 2713
rect 8894 2679 8937 2713
rect 8817 2634 8937 2679
rect 8817 2600 8860 2634
rect 8894 2600 8937 2634
rect 8255 1470 8298 1504
rect 8332 1470 8375 1504
rect 8255 1430 8375 1470
rect 8255 1396 8298 1430
rect 8332 1396 8375 1430
rect 8255 1250 8375 1396
rect 8255 1144 8262 1250
rect 8368 1144 8375 1250
rect 8817 1504 8937 2600
rect 9002 4098 9182 4099
rect 9002 4064 9003 4098
rect 9037 4082 9075 4098
rect 9037 4064 9039 4082
rect 9002 4048 9039 4064
rect 9073 4064 9075 4082
rect 9109 4082 9147 4098
rect 9109 4064 9111 4082
rect 9073 4048 9111 4064
rect 9145 4064 9147 4082
rect 9181 4064 9182 4098
rect 9145 4048 9182 4064
rect 9002 4025 9182 4048
rect 9002 3991 9003 4025
rect 9037 4014 9075 4025
rect 9037 3991 9039 4014
rect 9002 3980 9039 3991
rect 9073 3991 9075 4014
rect 9109 4014 9147 4025
rect 9109 3991 9111 4014
rect 9073 3980 9111 3991
rect 9145 3991 9147 4014
rect 9181 3991 9182 4025
rect 9145 3980 9182 3991
rect 9002 3952 9182 3980
rect 9002 3918 9003 3952
rect 9037 3946 9075 3952
rect 9037 3918 9039 3946
rect 9002 3912 9039 3918
rect 9073 3918 9075 3946
rect 9109 3946 9147 3952
rect 9109 3918 9111 3946
rect 9073 3912 9111 3918
rect 9145 3918 9147 3946
rect 9181 3918 9182 3952
rect 9145 3912 9182 3918
rect 9002 3879 9182 3912
rect 9002 3845 9003 3879
rect 9037 3878 9075 3879
rect 9037 3845 9039 3878
rect 9002 3844 9039 3845
rect 9073 3845 9075 3878
rect 9109 3878 9147 3879
rect 9109 3845 9111 3878
rect 9073 3844 9111 3845
rect 9145 3845 9147 3878
rect 9181 3845 9182 3879
rect 9145 3844 9182 3845
rect 9002 3810 9182 3844
rect 9002 3806 9039 3810
rect 9002 3772 9003 3806
rect 9037 3776 9039 3806
rect 9073 3806 9111 3810
rect 9073 3776 9075 3806
rect 9037 3772 9075 3776
rect 9109 3776 9111 3806
rect 9145 3806 9182 3810
rect 9145 3776 9147 3806
rect 9109 3772 9147 3776
rect 9181 3772 9182 3806
rect 9002 3742 9182 3772
rect 9002 3733 9039 3742
rect 9002 3699 9003 3733
rect 9037 3708 9039 3733
rect 9073 3733 9111 3742
rect 9073 3708 9075 3733
rect 9037 3699 9075 3708
rect 9109 3708 9111 3733
rect 9145 3733 9182 3742
rect 9145 3708 9147 3733
rect 9109 3699 9147 3708
rect 9181 3699 9182 3733
rect 9002 3674 9182 3699
rect 9002 3660 9039 3674
rect 9002 3626 9003 3660
rect 9037 3640 9039 3660
rect 9073 3660 9111 3674
rect 9073 3640 9075 3660
rect 9037 3626 9075 3640
rect 9109 3640 9111 3660
rect 9145 3660 9182 3674
rect 9145 3640 9147 3660
rect 9109 3626 9147 3640
rect 9181 3626 9182 3660
rect 9002 3606 9182 3626
rect 9002 3587 9039 3606
rect 9002 3553 9003 3587
rect 9037 3572 9039 3587
rect 9073 3587 9111 3606
rect 9073 3572 9075 3587
rect 9037 3553 9075 3572
rect 9109 3572 9111 3587
rect 9145 3587 9182 3606
rect 9145 3572 9147 3587
rect 9109 3553 9147 3572
rect 9181 3553 9182 3587
rect 9002 3538 9182 3553
rect 9002 3514 9039 3538
rect 9002 3480 9003 3514
rect 9037 3504 9039 3514
rect 9073 3514 9111 3538
rect 9073 3504 9075 3514
rect 9037 3480 9075 3504
rect 9109 3504 9111 3514
rect 9145 3514 9182 3538
rect 9145 3504 9147 3514
rect 9109 3480 9147 3504
rect 9181 3480 9182 3514
rect 9002 3470 9182 3480
rect 9002 3441 9039 3470
rect 9002 3407 9003 3441
rect 9037 3436 9039 3441
rect 9073 3441 9111 3470
rect 9073 3436 9075 3441
rect 9037 3407 9075 3436
rect 9109 3436 9111 3441
rect 9145 3441 9182 3470
rect 9145 3436 9147 3441
rect 9109 3407 9147 3436
rect 9181 3407 9182 3441
rect 9002 3402 9182 3407
rect 9002 3368 9039 3402
rect 9073 3368 9111 3402
rect 9145 3368 9182 3402
rect 9002 3334 9003 3368
rect 9037 3334 9075 3368
rect 9109 3334 9147 3368
rect 9181 3334 9182 3368
rect 9002 3300 9039 3334
rect 9073 3300 9111 3334
rect 9145 3300 9182 3334
rect 9002 3295 9182 3300
rect 9002 3261 9003 3295
rect 9037 3266 9075 3295
rect 9037 3261 9039 3266
rect 9002 3232 9039 3261
rect 9073 3261 9075 3266
rect 9109 3266 9147 3295
rect 9109 3261 9111 3266
rect 9073 3232 9111 3261
rect 9145 3261 9147 3266
rect 9181 3261 9182 3295
rect 9145 3232 9182 3261
rect 9002 3222 9182 3232
rect 9002 3188 9003 3222
rect 9037 3198 9075 3222
rect 9037 3188 9039 3198
rect 9002 3164 9039 3188
rect 9073 3188 9075 3198
rect 9109 3198 9147 3222
rect 9109 3188 9111 3198
rect 9073 3164 9111 3188
rect 9145 3188 9147 3198
rect 9181 3188 9182 3222
rect 9145 3164 9182 3188
rect 9002 3149 9182 3164
rect 9002 3115 9003 3149
rect 9037 3115 9075 3149
rect 9109 3115 9147 3149
rect 9181 3115 9182 3149
rect 9002 3076 9182 3115
rect 9002 3042 9003 3076
rect 9037 3042 9075 3076
rect 9109 3042 9147 3076
rect 9181 3042 9182 3076
rect 9002 3003 9182 3042
rect 9002 2969 9003 3003
rect 9037 2969 9075 3003
rect 9109 2969 9147 3003
rect 9181 2969 9182 3003
rect 9002 2930 9182 2969
rect 9002 2896 9003 2930
rect 9037 2896 9075 2930
rect 9109 2896 9147 2930
rect 9181 2896 9182 2930
rect 9002 2857 9182 2896
rect 9002 2823 9003 2857
rect 9037 2823 9075 2857
rect 9109 2823 9147 2857
rect 9181 2823 9182 2857
rect 9002 2784 9182 2823
rect 9002 2750 9003 2784
rect 9037 2750 9075 2784
rect 9109 2750 9147 2784
rect 9181 2750 9182 2784
rect 9002 2711 9182 2750
rect 9002 2677 9003 2711
rect 9037 2677 9075 2711
rect 9109 2677 9147 2711
rect 9181 2677 9182 2711
rect 9002 2638 9182 2677
rect 9002 2604 9003 2638
rect 9037 2604 9075 2638
rect 9109 2604 9147 2638
rect 9181 2604 9182 2638
rect 9002 2565 9182 2604
rect 9002 2531 9003 2565
rect 9037 2531 9075 2565
rect 9109 2531 9147 2565
rect 9181 2531 9182 2565
rect 9002 2492 9182 2531
rect 9002 2458 9003 2492
rect 9037 2482 9075 2492
rect 9037 2458 9039 2482
rect 9002 2448 9039 2458
rect 9073 2458 9075 2482
rect 9109 2482 9147 2492
rect 9109 2458 9111 2482
rect 9073 2448 9111 2458
rect 9145 2458 9147 2482
rect 9181 2458 9182 2492
rect 9145 2448 9182 2458
rect 9002 2419 9182 2448
rect 9002 2385 9003 2419
rect 9037 2414 9075 2419
rect 9037 2385 9039 2414
rect 9002 2380 9039 2385
rect 9073 2385 9075 2414
rect 9109 2414 9147 2419
rect 9109 2385 9111 2414
rect 9073 2380 9111 2385
rect 9145 2385 9147 2414
rect 9181 2385 9182 2419
rect 9145 2380 9182 2385
rect 9002 2346 9182 2380
rect 9002 2312 9003 2346
rect 9037 2312 9039 2346
rect 9073 2312 9075 2346
rect 9109 2312 9111 2346
rect 9145 2312 9147 2346
rect 9181 2312 9182 2346
rect 9002 2278 9182 2312
rect 9002 2273 9039 2278
rect 9002 2239 9003 2273
rect 9037 2244 9039 2273
rect 9073 2273 9111 2278
rect 9073 2244 9075 2273
rect 9037 2239 9075 2244
rect 9109 2244 9111 2273
rect 9145 2273 9182 2278
rect 9145 2244 9147 2273
rect 9109 2239 9147 2244
rect 9181 2239 9182 2273
rect 9002 2210 9182 2239
rect 9002 2200 9039 2210
rect 9002 2166 9003 2200
rect 9037 2176 9039 2200
rect 9073 2200 9111 2210
rect 9073 2176 9075 2200
rect 9037 2166 9075 2176
rect 9109 2176 9111 2200
rect 9145 2200 9182 2210
rect 9145 2176 9147 2200
rect 9109 2166 9147 2176
rect 9181 2166 9182 2200
rect 9002 2142 9182 2166
rect 9002 2126 9039 2142
rect 9002 2092 9003 2126
rect 9037 2108 9039 2126
rect 9073 2126 9111 2142
rect 9073 2108 9075 2126
rect 9037 2092 9075 2108
rect 9109 2108 9111 2126
rect 9145 2126 9182 2142
rect 9145 2108 9147 2126
rect 9109 2092 9147 2108
rect 9181 2092 9182 2126
rect 9002 2074 9182 2092
rect 9002 2052 9039 2074
rect 9002 2018 9003 2052
rect 9037 2040 9039 2052
rect 9073 2052 9111 2074
rect 9073 2040 9075 2052
rect 9037 2018 9075 2040
rect 9109 2040 9111 2052
rect 9145 2052 9182 2074
rect 9145 2040 9147 2052
rect 9109 2018 9147 2040
rect 9181 2018 9182 2052
rect 9002 2006 9182 2018
rect 9002 1978 9039 2006
rect 9002 1944 9003 1978
rect 9037 1972 9039 1978
rect 9073 1978 9111 2006
rect 9073 1972 9075 1978
rect 9037 1944 9075 1972
rect 9109 1972 9111 1978
rect 9145 1978 9182 2006
rect 9145 1972 9147 1978
rect 9109 1944 9147 1972
rect 9181 1944 9182 1978
rect 9002 1938 9182 1944
rect 9002 1904 9039 1938
rect 9073 1904 9111 1938
rect 9145 1904 9182 1938
rect 9002 1870 9003 1904
rect 9037 1870 9075 1904
rect 9109 1870 9147 1904
rect 9181 1870 9182 1904
rect 9002 1836 9039 1870
rect 9073 1836 9111 1870
rect 9145 1836 9182 1870
rect 9002 1830 9182 1836
rect 9002 1796 9003 1830
rect 9037 1802 9075 1830
rect 9037 1796 9039 1802
rect 9002 1768 9039 1796
rect 9073 1796 9075 1802
rect 9109 1802 9147 1830
rect 9109 1796 9111 1802
rect 9073 1768 9111 1796
rect 9145 1796 9147 1802
rect 9181 1796 9182 1830
rect 9145 1768 9182 1796
rect 9002 1756 9182 1768
rect 9002 1722 9003 1756
rect 9037 1734 9075 1756
rect 9037 1722 9039 1734
rect 9002 1700 9039 1722
rect 9073 1722 9075 1734
rect 9109 1734 9147 1756
rect 9109 1722 9111 1734
rect 9073 1700 9111 1722
rect 9145 1722 9147 1734
rect 9181 1722 9182 1756
rect 9145 1700 9182 1722
rect 9002 1682 9182 1700
rect 9002 1648 9003 1682
rect 9037 1666 9075 1682
rect 9037 1648 9039 1666
rect 9002 1632 9039 1648
rect 9073 1648 9075 1666
rect 9109 1666 9147 1682
rect 9109 1648 9111 1666
rect 9073 1632 9111 1648
rect 9145 1648 9147 1666
rect 9181 1648 9182 1682
rect 9145 1632 9182 1648
rect 9002 1608 9182 1632
rect 9002 1574 9003 1608
rect 9037 1598 9075 1608
rect 9037 1574 9039 1598
rect 9002 1564 9039 1574
rect 9073 1574 9075 1598
rect 9109 1598 9147 1608
rect 9109 1574 9111 1598
rect 9073 1564 9111 1574
rect 9145 1574 9147 1598
rect 9181 1574 9182 1608
rect 9145 1564 9182 1574
rect 9002 1548 9182 1564
rect 9247 3104 9367 4200
rect 9809 4308 9929 4324
rect 9809 4274 9852 4308
rect 9886 4274 9929 4308
rect 9809 4234 9929 4274
rect 9809 4200 9852 4234
rect 9886 4200 9929 4234
rect 9247 3070 9290 3104
rect 9324 3070 9367 3104
rect 9247 3026 9367 3070
rect 9247 2992 9290 3026
rect 9324 2992 9367 3026
rect 9247 2948 9367 2992
rect 9247 2914 9290 2948
rect 9324 2914 9367 2948
rect 9247 2870 9367 2914
rect 9247 2836 9290 2870
rect 9324 2836 9367 2870
rect 9247 2792 9367 2836
rect 9247 2758 9290 2792
rect 9324 2758 9367 2792
rect 9247 2713 9367 2758
rect 9247 2679 9290 2713
rect 9324 2679 9367 2713
rect 9247 2634 9367 2679
rect 9247 2600 9290 2634
rect 9324 2600 9367 2634
rect 8817 1470 8860 1504
rect 8894 1470 8937 1504
rect 8817 1430 8937 1470
rect 8817 1396 8860 1430
rect 8894 1396 8937 1430
rect 8817 1250 8937 1396
rect 8817 1144 8824 1250
rect 8930 1144 8937 1250
rect 9247 1504 9367 2600
rect 9469 4092 9571 4118
rect 9605 4092 9707 4118
rect 9469 4082 9499 4092
rect 9677 4082 9707 4092
rect 9469 4014 9499 4048
rect 9677 4014 9707 4048
rect 9469 3946 9499 3980
rect 9677 3946 9707 3980
rect 9469 3878 9499 3912
rect 9677 3878 9707 3912
rect 9469 3810 9499 3844
rect 9677 3810 9707 3844
rect 9469 3742 9499 3776
rect 9677 3742 9707 3776
rect 9469 3674 9499 3708
rect 9677 3674 9707 3708
rect 9469 3606 9499 3640
rect 9677 3606 9707 3640
rect 9469 3538 9499 3572
rect 9677 3538 9707 3572
rect 9469 3470 9499 3504
rect 9677 3470 9707 3504
rect 9469 3402 9499 3436
rect 9677 3402 9707 3436
rect 9469 3334 9499 3368
rect 9677 3334 9707 3368
rect 9469 3266 9499 3300
rect 9677 3266 9707 3300
rect 9469 3198 9499 3232
rect 9677 3198 9707 3232
rect 9503 3164 9571 3194
rect 9605 3164 9673 3194
rect 9469 3148 9571 3164
rect 9605 3148 9707 3164
rect 9469 3108 9707 3148
rect 9469 3074 9499 3108
rect 9533 3074 9571 3108
rect 9605 3074 9643 3108
rect 9677 3074 9707 3108
rect 9469 3044 9707 3074
rect 9469 3028 9537 3044
rect 9469 2994 9499 3028
rect 9533 3010 9537 3028
rect 9571 3028 9605 3044
rect 9533 2994 9571 3010
rect 9639 3028 9707 3044
rect 9639 3010 9643 3028
rect 9605 2994 9643 3010
rect 9677 2994 9707 3028
rect 9469 2974 9707 2994
rect 9469 2948 9537 2974
rect 9469 2914 9499 2948
rect 9533 2940 9537 2948
rect 9571 2948 9605 2974
rect 9533 2914 9571 2940
rect 9639 2948 9707 2974
rect 9639 2940 9643 2948
rect 9605 2914 9643 2940
rect 9677 2914 9707 2948
rect 9469 2904 9707 2914
rect 9469 2870 9537 2904
rect 9571 2870 9605 2904
rect 9639 2870 9707 2904
rect 9469 2868 9707 2870
rect 9469 2834 9499 2868
rect 9533 2834 9571 2868
rect 9605 2834 9643 2868
rect 9677 2834 9707 2868
rect 9469 2800 9537 2834
rect 9571 2800 9605 2834
rect 9639 2800 9707 2834
rect 9469 2788 9707 2800
rect 9469 2754 9499 2788
rect 9533 2764 9571 2788
rect 9533 2754 9537 2764
rect 9469 2730 9537 2754
rect 9605 2764 9643 2788
rect 9571 2730 9605 2754
rect 9639 2754 9643 2764
rect 9677 2754 9707 2788
rect 9639 2730 9707 2754
rect 9469 2708 9707 2730
rect 9469 2674 9499 2708
rect 9533 2694 9571 2708
rect 9533 2674 9537 2694
rect 9469 2660 9537 2674
rect 9605 2694 9643 2708
rect 9571 2660 9605 2674
rect 9639 2674 9643 2694
rect 9677 2674 9707 2708
rect 9639 2660 9707 2674
rect 9469 2628 9707 2660
rect 9469 2594 9499 2628
rect 9533 2594 9571 2628
rect 9605 2594 9643 2628
rect 9677 2594 9707 2628
rect 9469 2556 9707 2594
rect 9469 2540 9571 2556
rect 9605 2540 9707 2556
rect 9503 2518 9571 2540
rect 9605 2518 9673 2540
rect 9469 2472 9499 2506
rect 9677 2472 9707 2506
rect 9469 2404 9499 2438
rect 9677 2404 9707 2438
rect 9469 2336 9499 2370
rect 9677 2336 9707 2370
rect 9469 2268 9499 2302
rect 9677 2268 9707 2302
rect 9469 2200 9499 2234
rect 9677 2200 9707 2234
rect 9469 2132 9499 2166
rect 9677 2132 9707 2166
rect 9469 2064 9499 2098
rect 9677 2064 9707 2098
rect 9469 1996 9499 2030
rect 9677 1996 9707 2030
rect 9469 1928 9499 1962
rect 9677 1928 9707 1962
rect 9469 1860 9499 1894
rect 9677 1860 9707 1894
rect 9469 1792 9499 1826
rect 9677 1792 9707 1826
rect 9469 1724 9499 1758
rect 9677 1724 9707 1758
rect 9469 1656 9499 1690
rect 9677 1656 9707 1690
rect 9469 1620 9499 1622
rect 9677 1620 9707 1622
rect 9469 1586 9571 1620
rect 9605 1586 9707 1620
rect 9469 1536 9707 1586
rect 9809 3104 9929 4200
rect 10239 4308 10359 4324
rect 10239 4274 10282 4308
rect 10316 4274 10359 4308
rect 10239 4234 10359 4274
rect 10239 4200 10282 4234
rect 10316 4200 10359 4234
rect 9809 3070 9852 3104
rect 9886 3070 9929 3104
rect 9809 3026 9929 3070
rect 9809 2992 9852 3026
rect 9886 2992 9929 3026
rect 9809 2948 9929 2992
rect 9809 2914 9852 2948
rect 9886 2914 9929 2948
rect 9809 2870 9929 2914
rect 9809 2836 9852 2870
rect 9886 2836 9929 2870
rect 9809 2792 9929 2836
rect 9809 2758 9852 2792
rect 9886 2758 9929 2792
rect 9809 2713 9929 2758
rect 9809 2679 9852 2713
rect 9886 2679 9929 2713
rect 9809 2634 9929 2679
rect 9809 2600 9852 2634
rect 9886 2600 9929 2634
rect 9247 1470 9290 1504
rect 9324 1470 9367 1504
rect 9247 1430 9367 1470
rect 9247 1396 9290 1430
rect 9324 1396 9367 1430
rect 9247 1250 9367 1396
rect 9247 1144 9254 1250
rect 9360 1144 9367 1250
rect 9809 1504 9929 2600
rect 9994 4098 10174 4118
rect 9994 4064 9995 4098
rect 10029 4082 10067 4098
rect 10029 4064 10031 4082
rect 9994 4048 10031 4064
rect 10065 4064 10067 4082
rect 10101 4082 10139 4098
rect 10101 4064 10103 4082
rect 10065 4048 10103 4064
rect 10137 4064 10139 4082
rect 10173 4064 10174 4098
rect 10137 4048 10174 4064
rect 9994 4025 10174 4048
rect 9994 3991 9995 4025
rect 10029 4014 10067 4025
rect 10029 3991 10031 4014
rect 9994 3980 10031 3991
rect 10065 3991 10067 4014
rect 10101 4014 10139 4025
rect 10101 3991 10103 4014
rect 10065 3980 10103 3991
rect 10137 3991 10139 4014
rect 10173 3991 10174 4025
rect 10137 3980 10174 3991
rect 9994 3952 10174 3980
rect 9994 3918 9995 3952
rect 10029 3946 10067 3952
rect 10029 3918 10031 3946
rect 9994 3912 10031 3918
rect 10065 3918 10067 3946
rect 10101 3946 10139 3952
rect 10101 3918 10103 3946
rect 10065 3912 10103 3918
rect 10137 3918 10139 3946
rect 10173 3918 10174 3952
rect 10137 3912 10174 3918
rect 9994 3879 10174 3912
rect 9994 3845 9995 3879
rect 10029 3878 10067 3879
rect 10029 3845 10031 3878
rect 9994 3844 10031 3845
rect 10065 3845 10067 3878
rect 10101 3878 10139 3879
rect 10101 3845 10103 3878
rect 10065 3844 10103 3845
rect 10137 3845 10139 3878
rect 10173 3845 10174 3879
rect 10137 3844 10174 3845
rect 9994 3810 10174 3844
rect 9994 3806 10031 3810
rect 9994 3772 9995 3806
rect 10029 3776 10031 3806
rect 10065 3806 10103 3810
rect 10065 3776 10067 3806
rect 10029 3772 10067 3776
rect 10101 3776 10103 3806
rect 10137 3806 10174 3810
rect 10137 3776 10139 3806
rect 10101 3772 10139 3776
rect 10173 3772 10174 3806
rect 9994 3742 10174 3772
rect 9994 3733 10031 3742
rect 9994 3699 9995 3733
rect 10029 3708 10031 3733
rect 10065 3733 10103 3742
rect 10065 3708 10067 3733
rect 10029 3699 10067 3708
rect 10101 3708 10103 3733
rect 10137 3733 10174 3742
rect 10137 3708 10139 3733
rect 10101 3699 10139 3708
rect 10173 3699 10174 3733
rect 9994 3674 10174 3699
rect 9994 3660 10031 3674
rect 9994 3626 9995 3660
rect 10029 3640 10031 3660
rect 10065 3660 10103 3674
rect 10065 3640 10067 3660
rect 10029 3626 10067 3640
rect 10101 3640 10103 3660
rect 10137 3660 10174 3674
rect 10137 3640 10139 3660
rect 10101 3626 10139 3640
rect 10173 3626 10174 3660
rect 9994 3606 10174 3626
rect 9994 3587 10031 3606
rect 9994 3553 9995 3587
rect 10029 3572 10031 3587
rect 10065 3587 10103 3606
rect 10065 3572 10067 3587
rect 10029 3553 10067 3572
rect 10101 3572 10103 3587
rect 10137 3587 10174 3606
rect 10137 3572 10139 3587
rect 10101 3553 10139 3572
rect 10173 3553 10174 3587
rect 9994 3538 10174 3553
rect 9994 3514 10031 3538
rect 9994 3480 9995 3514
rect 10029 3504 10031 3514
rect 10065 3514 10103 3538
rect 10065 3504 10067 3514
rect 10029 3480 10067 3504
rect 10101 3504 10103 3514
rect 10137 3514 10174 3538
rect 10137 3504 10139 3514
rect 10101 3480 10139 3504
rect 10173 3480 10174 3514
rect 9994 3470 10174 3480
rect 9994 3441 10031 3470
rect 9994 3407 9995 3441
rect 10029 3436 10031 3441
rect 10065 3441 10103 3470
rect 10065 3436 10067 3441
rect 10029 3407 10067 3436
rect 10101 3436 10103 3441
rect 10137 3441 10174 3470
rect 10137 3436 10139 3441
rect 10101 3407 10139 3436
rect 10173 3407 10174 3441
rect 9994 3402 10174 3407
rect 9994 3368 10031 3402
rect 10065 3368 10103 3402
rect 10137 3368 10174 3402
rect 9994 3334 9995 3368
rect 10029 3334 10067 3368
rect 10101 3334 10139 3368
rect 10173 3334 10174 3368
rect 9994 3300 10031 3334
rect 10065 3300 10103 3334
rect 10137 3300 10174 3334
rect 9994 3295 10174 3300
rect 9994 3261 9995 3295
rect 10029 3266 10067 3295
rect 10029 3261 10031 3266
rect 9994 3232 10031 3261
rect 10065 3261 10067 3266
rect 10101 3266 10139 3295
rect 10101 3261 10103 3266
rect 10065 3232 10103 3261
rect 10137 3261 10139 3266
rect 10173 3261 10174 3295
rect 10137 3232 10174 3261
rect 9994 3222 10174 3232
rect 9994 3188 9995 3222
rect 10029 3198 10067 3222
rect 10029 3188 10031 3198
rect 9994 3164 10031 3188
rect 10065 3188 10067 3198
rect 10101 3198 10139 3222
rect 10101 3188 10103 3198
rect 10065 3164 10103 3188
rect 10137 3188 10139 3198
rect 10173 3188 10174 3222
rect 10137 3164 10174 3188
rect 9994 3149 10174 3164
rect 9994 3115 9995 3149
rect 10029 3115 10067 3149
rect 10101 3115 10139 3149
rect 10173 3115 10174 3149
rect 9994 3076 10174 3115
rect 9994 3042 9995 3076
rect 10029 3042 10067 3076
rect 10101 3042 10139 3076
rect 10173 3042 10174 3076
rect 9994 3003 10174 3042
rect 9994 2969 9995 3003
rect 10029 2969 10067 3003
rect 10101 2969 10139 3003
rect 10173 2969 10174 3003
rect 9994 2930 10174 2969
rect 9994 2896 9995 2930
rect 10029 2896 10067 2930
rect 10101 2896 10139 2930
rect 10173 2896 10174 2930
rect 9994 2857 10174 2896
rect 9994 2823 9995 2857
rect 10029 2823 10067 2857
rect 10101 2823 10139 2857
rect 10173 2823 10174 2857
rect 9994 2784 10174 2823
rect 9994 2750 9995 2784
rect 10029 2750 10067 2784
rect 10101 2750 10139 2784
rect 10173 2750 10174 2784
rect 9994 2711 10174 2750
rect 9994 2677 9995 2711
rect 10029 2677 10067 2711
rect 10101 2677 10139 2711
rect 10173 2677 10174 2711
rect 9994 2638 10174 2677
rect 9994 2604 9995 2638
rect 10029 2604 10067 2638
rect 10101 2604 10139 2638
rect 10173 2604 10174 2638
rect 9994 2565 10174 2604
rect 9994 2531 9995 2565
rect 10029 2531 10067 2565
rect 10101 2531 10139 2565
rect 10173 2531 10174 2565
rect 9994 2492 10174 2531
rect 9994 2458 9995 2492
rect 10029 2482 10067 2492
rect 10029 2458 10031 2482
rect 9994 2448 10031 2458
rect 10065 2458 10067 2482
rect 10101 2482 10139 2492
rect 10101 2458 10103 2482
rect 10065 2448 10103 2458
rect 10137 2458 10139 2482
rect 10173 2458 10174 2492
rect 10137 2448 10174 2458
rect 9994 2419 10174 2448
rect 9994 2385 9995 2419
rect 10029 2414 10067 2419
rect 10029 2385 10031 2414
rect 9994 2380 10031 2385
rect 10065 2385 10067 2414
rect 10101 2414 10139 2419
rect 10101 2385 10103 2414
rect 10065 2380 10103 2385
rect 10137 2385 10139 2414
rect 10173 2385 10174 2419
rect 10137 2380 10174 2385
rect 9994 2346 10174 2380
rect 9994 2312 9995 2346
rect 10029 2312 10031 2346
rect 10065 2312 10067 2346
rect 10101 2312 10103 2346
rect 10137 2312 10139 2346
rect 10173 2312 10174 2346
rect 9994 2278 10174 2312
rect 9994 2273 10031 2278
rect 9994 2239 9995 2273
rect 10029 2244 10031 2273
rect 10065 2273 10103 2278
rect 10065 2244 10067 2273
rect 10029 2239 10067 2244
rect 10101 2244 10103 2273
rect 10137 2273 10174 2278
rect 10137 2244 10139 2273
rect 10101 2239 10139 2244
rect 10173 2239 10174 2273
rect 9994 2210 10174 2239
rect 9994 2200 10031 2210
rect 9994 2166 9995 2200
rect 10029 2176 10031 2200
rect 10065 2200 10103 2210
rect 10065 2176 10067 2200
rect 10029 2166 10067 2176
rect 10101 2176 10103 2200
rect 10137 2200 10174 2210
rect 10137 2176 10139 2200
rect 10101 2166 10139 2176
rect 10173 2166 10174 2200
rect 9994 2142 10174 2166
rect 9994 2126 10031 2142
rect 9994 2092 9995 2126
rect 10029 2108 10031 2126
rect 10065 2126 10103 2142
rect 10065 2108 10067 2126
rect 10029 2092 10067 2108
rect 10101 2108 10103 2126
rect 10137 2126 10174 2142
rect 10137 2108 10139 2126
rect 10101 2092 10139 2108
rect 10173 2092 10174 2126
rect 9994 2074 10174 2092
rect 9994 2052 10031 2074
rect 9994 2018 9995 2052
rect 10029 2040 10031 2052
rect 10065 2052 10103 2074
rect 10065 2040 10067 2052
rect 10029 2018 10067 2040
rect 10101 2040 10103 2052
rect 10137 2052 10174 2074
rect 10137 2040 10139 2052
rect 10101 2018 10139 2040
rect 10173 2018 10174 2052
rect 9994 2006 10174 2018
rect 9994 1978 10031 2006
rect 9994 1944 9995 1978
rect 10029 1972 10031 1978
rect 10065 1978 10103 2006
rect 10065 1972 10067 1978
rect 10029 1944 10067 1972
rect 10101 1972 10103 1978
rect 10137 1978 10174 2006
rect 10137 1972 10139 1978
rect 10101 1944 10139 1972
rect 10173 1944 10174 1978
rect 9994 1938 10174 1944
rect 9994 1904 10031 1938
rect 10065 1904 10103 1938
rect 10137 1904 10174 1938
rect 9994 1870 9995 1904
rect 10029 1870 10067 1904
rect 10101 1870 10139 1904
rect 10173 1870 10174 1904
rect 9994 1836 10031 1870
rect 10065 1836 10103 1870
rect 10137 1836 10174 1870
rect 9994 1830 10174 1836
rect 9994 1796 9995 1830
rect 10029 1802 10067 1830
rect 10029 1796 10031 1802
rect 9994 1768 10031 1796
rect 10065 1796 10067 1802
rect 10101 1802 10139 1830
rect 10101 1796 10103 1802
rect 10065 1768 10103 1796
rect 10137 1796 10139 1802
rect 10173 1796 10174 1830
rect 10137 1768 10174 1796
rect 9994 1756 10174 1768
rect 9994 1722 9995 1756
rect 10029 1734 10067 1756
rect 10029 1722 10031 1734
rect 9994 1700 10031 1722
rect 10065 1722 10067 1734
rect 10101 1734 10139 1756
rect 10101 1722 10103 1734
rect 10065 1700 10103 1722
rect 10137 1722 10139 1734
rect 10173 1722 10174 1756
rect 10137 1700 10174 1722
rect 9994 1682 10174 1700
rect 9994 1648 9995 1682
rect 10029 1666 10067 1682
rect 10029 1648 10031 1666
rect 9994 1632 10031 1648
rect 10065 1648 10067 1666
rect 10101 1666 10139 1682
rect 10101 1648 10103 1666
rect 10065 1632 10103 1648
rect 10137 1648 10139 1666
rect 10173 1648 10174 1682
rect 10137 1632 10174 1648
rect 9994 1608 10174 1632
rect 9994 1574 9995 1608
rect 10029 1598 10067 1608
rect 10029 1574 10031 1598
rect 9994 1564 10031 1574
rect 10065 1574 10067 1598
rect 10101 1598 10139 1608
rect 10101 1574 10103 1598
rect 10065 1564 10103 1574
rect 10137 1574 10139 1598
rect 10173 1574 10174 1608
rect 10137 1564 10174 1574
rect 9994 1548 10174 1564
rect 10239 3104 10359 4200
rect 10801 4308 10921 4324
rect 10801 4274 10844 4308
rect 10878 4274 10921 4308
rect 10801 4234 10921 4274
rect 10801 4200 10844 4234
rect 10878 4200 10921 4234
rect 10239 3070 10282 3104
rect 10316 3070 10359 3104
rect 10239 3026 10359 3070
rect 10239 2992 10282 3026
rect 10316 2992 10359 3026
rect 10239 2948 10359 2992
rect 10239 2914 10282 2948
rect 10316 2914 10359 2948
rect 10239 2870 10359 2914
rect 10239 2836 10282 2870
rect 10316 2836 10359 2870
rect 10239 2792 10359 2836
rect 10239 2758 10282 2792
rect 10316 2758 10359 2792
rect 10239 2713 10359 2758
rect 10239 2679 10282 2713
rect 10316 2679 10359 2713
rect 10239 2634 10359 2679
rect 10239 2600 10282 2634
rect 10316 2600 10359 2634
rect 9809 1470 9852 1504
rect 9886 1470 9929 1504
rect 9809 1430 9929 1470
rect 9809 1396 9852 1430
rect 9886 1396 9929 1430
rect 9809 1250 9929 1396
rect 9809 1144 9816 1250
rect 9922 1144 9929 1250
rect 10239 1504 10359 2600
rect 10461 4118 10699 4130
rect 10461 4092 10563 4118
rect 10597 4092 10699 4118
rect 10461 4082 10491 4092
rect 10669 4082 10699 4092
rect 10461 4014 10491 4048
rect 10669 4014 10699 4048
rect 10461 3946 10491 3980
rect 10669 3946 10699 3980
rect 10461 3878 10491 3912
rect 10669 3878 10699 3912
rect 10461 3810 10491 3844
rect 10669 3810 10699 3844
rect 10461 3742 10491 3776
rect 10669 3742 10699 3776
rect 10461 3674 10491 3708
rect 10669 3674 10699 3708
rect 10461 3606 10491 3640
rect 10669 3606 10699 3640
rect 10461 3538 10491 3572
rect 10669 3538 10699 3572
rect 10461 3470 10491 3504
rect 10669 3470 10699 3504
rect 10461 3402 10491 3436
rect 10669 3402 10699 3436
rect 10461 3334 10491 3368
rect 10669 3334 10699 3368
rect 10461 3266 10491 3300
rect 10669 3266 10699 3300
rect 10461 3198 10491 3232
rect 10669 3198 10699 3232
rect 10495 3164 10563 3194
rect 10597 3164 10665 3194
rect 10461 3148 10563 3164
rect 10597 3148 10699 3164
rect 10461 3108 10699 3148
rect 10461 3074 10491 3108
rect 10525 3074 10563 3108
rect 10597 3074 10635 3108
rect 10669 3074 10699 3108
rect 10461 3044 10699 3074
rect 10461 3028 10529 3044
rect 10461 2994 10491 3028
rect 10525 3010 10529 3028
rect 10563 3028 10597 3044
rect 10525 2994 10563 3010
rect 10631 3028 10699 3044
rect 10631 3010 10635 3028
rect 10597 2994 10635 3010
rect 10669 2994 10699 3028
rect 10461 2974 10699 2994
rect 10461 2948 10529 2974
rect 10461 2914 10491 2948
rect 10525 2940 10529 2948
rect 10563 2948 10597 2974
rect 10525 2914 10563 2940
rect 10631 2948 10699 2974
rect 10631 2940 10635 2948
rect 10597 2914 10635 2940
rect 10669 2914 10699 2948
rect 10461 2904 10699 2914
rect 10461 2870 10529 2904
rect 10563 2870 10597 2904
rect 10631 2870 10699 2904
rect 10461 2868 10699 2870
rect 10461 2834 10491 2868
rect 10525 2834 10563 2868
rect 10597 2834 10635 2868
rect 10669 2834 10699 2868
rect 10461 2800 10529 2834
rect 10563 2800 10597 2834
rect 10631 2800 10699 2834
rect 10461 2788 10699 2800
rect 10461 2754 10491 2788
rect 10525 2764 10563 2788
rect 10525 2754 10529 2764
rect 10461 2730 10529 2754
rect 10597 2764 10635 2788
rect 10563 2730 10597 2754
rect 10631 2754 10635 2764
rect 10669 2754 10699 2788
rect 10631 2730 10699 2754
rect 10461 2708 10699 2730
rect 10461 2674 10491 2708
rect 10525 2694 10563 2708
rect 10525 2674 10529 2694
rect 10461 2660 10529 2674
rect 10597 2694 10635 2708
rect 10563 2660 10597 2674
rect 10631 2674 10635 2694
rect 10669 2674 10699 2708
rect 10631 2660 10699 2674
rect 10461 2628 10699 2660
rect 10461 2594 10491 2628
rect 10525 2594 10563 2628
rect 10597 2594 10635 2628
rect 10669 2594 10699 2628
rect 10461 2556 10699 2594
rect 10461 2540 10563 2556
rect 10597 2540 10699 2556
rect 10495 2518 10563 2540
rect 10597 2518 10665 2540
rect 10461 2472 10491 2506
rect 10669 2472 10699 2506
rect 10461 2404 10491 2438
rect 10669 2404 10699 2438
rect 10461 2336 10491 2370
rect 10669 2336 10699 2370
rect 10461 2268 10491 2302
rect 10669 2268 10699 2302
rect 10461 2200 10491 2234
rect 10669 2200 10699 2234
rect 10461 2132 10491 2166
rect 10669 2132 10699 2166
rect 10461 2064 10491 2098
rect 10669 2064 10699 2098
rect 10461 1996 10491 2030
rect 10669 1996 10699 2030
rect 10461 1928 10491 1962
rect 10669 1928 10699 1962
rect 10461 1860 10491 1894
rect 10669 1860 10699 1894
rect 10461 1792 10491 1826
rect 10669 1792 10699 1826
rect 10461 1724 10491 1758
rect 10669 1724 10699 1758
rect 10461 1656 10491 1690
rect 10669 1656 10699 1690
rect 10461 1620 10491 1622
rect 10669 1620 10699 1622
rect 10461 1586 10563 1620
rect 10597 1586 10699 1620
rect 10461 1536 10699 1586
rect 10801 3104 10921 4200
rect 11231 4308 11351 4324
rect 11231 4274 11274 4308
rect 11308 4274 11351 4308
rect 11231 4234 11351 4274
rect 11231 4200 11274 4234
rect 11308 4200 11351 4234
rect 10801 3070 10844 3104
rect 10878 3070 10921 3104
rect 10801 3026 10921 3070
rect 10801 2992 10844 3026
rect 10878 2992 10921 3026
rect 10801 2948 10921 2992
rect 10801 2914 10844 2948
rect 10878 2914 10921 2948
rect 10801 2870 10921 2914
rect 10801 2836 10844 2870
rect 10878 2836 10921 2870
rect 10801 2792 10921 2836
rect 10801 2758 10844 2792
rect 10878 2758 10921 2792
rect 10801 2713 10921 2758
rect 10801 2679 10844 2713
rect 10878 2679 10921 2713
rect 10801 2634 10921 2679
rect 10801 2600 10844 2634
rect 10878 2600 10921 2634
rect 10239 1470 10282 1504
rect 10316 1470 10359 1504
rect 10239 1430 10359 1470
rect 10239 1396 10282 1430
rect 10316 1396 10359 1430
rect 10239 1250 10359 1396
rect 10239 1144 10246 1250
rect 10352 1144 10359 1250
rect 10801 1504 10921 2600
rect 10986 4064 10987 4098
rect 11021 4082 11059 4098
rect 11021 4064 11023 4082
rect 10986 4048 11023 4064
rect 11057 4064 11059 4082
rect 11093 4082 11131 4098
rect 11093 4064 11095 4082
rect 11057 4048 11095 4064
rect 11129 4064 11131 4082
rect 11165 4064 11166 4098
rect 11129 4048 11166 4064
rect 10986 4025 11166 4048
rect 10986 3991 10987 4025
rect 11021 4014 11059 4025
rect 11021 3991 11023 4014
rect 10986 3980 11023 3991
rect 11057 3991 11059 4014
rect 11093 4014 11131 4025
rect 11093 3991 11095 4014
rect 11057 3980 11095 3991
rect 11129 3991 11131 4014
rect 11165 3991 11166 4025
rect 11129 3980 11166 3991
rect 10986 3952 11166 3980
rect 10986 3918 10987 3952
rect 11021 3946 11059 3952
rect 11021 3918 11023 3946
rect 10986 3912 11023 3918
rect 11057 3918 11059 3946
rect 11093 3946 11131 3952
rect 11093 3918 11095 3946
rect 11057 3912 11095 3918
rect 11129 3918 11131 3946
rect 11165 3918 11166 3952
rect 11129 3912 11166 3918
rect 10986 3879 11166 3912
rect 10986 3845 10987 3879
rect 11021 3878 11059 3879
rect 11021 3845 11023 3878
rect 10986 3844 11023 3845
rect 11057 3845 11059 3878
rect 11093 3878 11131 3879
rect 11093 3845 11095 3878
rect 11057 3844 11095 3845
rect 11129 3845 11131 3878
rect 11165 3845 11166 3879
rect 11129 3844 11166 3845
rect 10986 3810 11166 3844
rect 10986 3806 11023 3810
rect 10986 3772 10987 3806
rect 11021 3776 11023 3806
rect 11057 3806 11095 3810
rect 11057 3776 11059 3806
rect 11021 3772 11059 3776
rect 11093 3776 11095 3806
rect 11129 3806 11166 3810
rect 11129 3776 11131 3806
rect 11093 3772 11131 3776
rect 11165 3772 11166 3806
rect 10986 3742 11166 3772
rect 10986 3733 11023 3742
rect 10986 3699 10987 3733
rect 11021 3708 11023 3733
rect 11057 3733 11095 3742
rect 11057 3708 11059 3733
rect 11021 3699 11059 3708
rect 11093 3708 11095 3733
rect 11129 3733 11166 3742
rect 11129 3708 11131 3733
rect 11093 3699 11131 3708
rect 11165 3699 11166 3733
rect 10986 3674 11166 3699
rect 10986 3660 11023 3674
rect 10986 3626 10987 3660
rect 11021 3640 11023 3660
rect 11057 3660 11095 3674
rect 11057 3640 11059 3660
rect 11021 3626 11059 3640
rect 11093 3640 11095 3660
rect 11129 3660 11166 3674
rect 11129 3640 11131 3660
rect 11093 3626 11131 3640
rect 11165 3626 11166 3660
rect 10986 3606 11166 3626
rect 10986 3587 11023 3606
rect 10986 3553 10987 3587
rect 11021 3572 11023 3587
rect 11057 3587 11095 3606
rect 11057 3572 11059 3587
rect 11021 3553 11059 3572
rect 11093 3572 11095 3587
rect 11129 3587 11166 3606
rect 11129 3572 11131 3587
rect 11093 3553 11131 3572
rect 11165 3553 11166 3587
rect 10986 3538 11166 3553
rect 10986 3514 11023 3538
rect 10986 3480 10987 3514
rect 11021 3504 11023 3514
rect 11057 3514 11095 3538
rect 11057 3504 11059 3514
rect 11021 3480 11059 3504
rect 11093 3504 11095 3514
rect 11129 3514 11166 3538
rect 11129 3504 11131 3514
rect 11093 3480 11131 3504
rect 11165 3480 11166 3514
rect 10986 3470 11166 3480
rect 10986 3441 11023 3470
rect 10986 3407 10987 3441
rect 11021 3436 11023 3441
rect 11057 3441 11095 3470
rect 11057 3436 11059 3441
rect 11021 3407 11059 3436
rect 11093 3436 11095 3441
rect 11129 3441 11166 3470
rect 11129 3436 11131 3441
rect 11093 3407 11131 3436
rect 11165 3407 11166 3441
rect 10986 3402 11166 3407
rect 10986 3368 11023 3402
rect 11057 3368 11095 3402
rect 11129 3368 11166 3402
rect 10986 3334 10987 3368
rect 11021 3334 11059 3368
rect 11093 3334 11131 3368
rect 11165 3334 11166 3368
rect 10986 3300 11023 3334
rect 11057 3300 11095 3334
rect 11129 3300 11166 3334
rect 10986 3295 11166 3300
rect 10986 3261 10987 3295
rect 11021 3266 11059 3295
rect 11021 3261 11023 3266
rect 10986 3232 11023 3261
rect 11057 3261 11059 3266
rect 11093 3266 11131 3295
rect 11093 3261 11095 3266
rect 11057 3232 11095 3261
rect 11129 3261 11131 3266
rect 11165 3261 11166 3295
rect 11129 3232 11166 3261
rect 10986 3222 11166 3232
rect 10986 3188 10987 3222
rect 11021 3198 11059 3222
rect 11021 3188 11023 3198
rect 10986 3164 11023 3188
rect 11057 3188 11059 3198
rect 11093 3198 11131 3222
rect 11093 3188 11095 3198
rect 11057 3164 11095 3188
rect 11129 3188 11131 3198
rect 11165 3188 11166 3222
rect 11129 3164 11166 3188
rect 10986 3149 11166 3164
rect 10986 3115 10987 3149
rect 11021 3115 11059 3149
rect 11093 3115 11131 3149
rect 11165 3115 11166 3149
rect 10986 3076 11166 3115
rect 10986 3042 10987 3076
rect 11021 3042 11059 3076
rect 11093 3042 11131 3076
rect 11165 3042 11166 3076
rect 10986 3003 11166 3042
rect 10986 2969 10987 3003
rect 11021 2969 11059 3003
rect 11093 2969 11131 3003
rect 11165 2969 11166 3003
rect 10986 2930 11166 2969
rect 10986 2896 10987 2930
rect 11021 2896 11059 2930
rect 11093 2896 11131 2930
rect 11165 2896 11166 2930
rect 10986 2857 11166 2896
rect 10986 2823 10987 2857
rect 11021 2823 11059 2857
rect 11093 2823 11131 2857
rect 11165 2823 11166 2857
rect 10986 2784 11166 2823
rect 10986 2750 10987 2784
rect 11021 2750 11059 2784
rect 11093 2750 11131 2784
rect 11165 2750 11166 2784
rect 10986 2711 11166 2750
rect 10986 2677 10987 2711
rect 11021 2677 11059 2711
rect 11093 2677 11131 2711
rect 11165 2677 11166 2711
rect 10986 2638 11166 2677
rect 10986 2604 10987 2638
rect 11021 2604 11059 2638
rect 11093 2604 11131 2638
rect 11165 2604 11166 2638
rect 10986 2565 11166 2604
rect 10986 2531 10987 2565
rect 11021 2531 11059 2565
rect 11093 2531 11131 2565
rect 11165 2531 11166 2565
rect 10986 2492 11166 2531
rect 10986 2458 10987 2492
rect 11021 2482 11059 2492
rect 11021 2458 11023 2482
rect 10986 2448 11023 2458
rect 11057 2458 11059 2482
rect 11093 2482 11131 2492
rect 11093 2458 11095 2482
rect 11057 2448 11095 2458
rect 11129 2458 11131 2482
rect 11165 2458 11166 2492
rect 11129 2448 11166 2458
rect 10986 2419 11166 2448
rect 10986 2385 10987 2419
rect 11021 2414 11059 2419
rect 11021 2385 11023 2414
rect 10986 2380 11023 2385
rect 11057 2385 11059 2414
rect 11093 2414 11131 2419
rect 11093 2385 11095 2414
rect 11057 2380 11095 2385
rect 11129 2385 11131 2414
rect 11165 2385 11166 2419
rect 11129 2380 11166 2385
rect 10986 2346 11166 2380
rect 10986 2312 10987 2346
rect 11021 2312 11023 2346
rect 11057 2312 11059 2346
rect 11093 2312 11095 2346
rect 11129 2312 11131 2346
rect 11165 2312 11166 2346
rect 10986 2278 11166 2312
rect 10986 2273 11023 2278
rect 10986 2239 10987 2273
rect 11021 2244 11023 2273
rect 11057 2273 11095 2278
rect 11057 2244 11059 2273
rect 11021 2239 11059 2244
rect 11093 2244 11095 2273
rect 11129 2273 11166 2278
rect 11129 2244 11131 2273
rect 11093 2239 11131 2244
rect 11165 2239 11166 2273
rect 10986 2210 11166 2239
rect 10986 2200 11023 2210
rect 10986 2166 10987 2200
rect 11021 2176 11023 2200
rect 11057 2200 11095 2210
rect 11057 2176 11059 2200
rect 11021 2166 11059 2176
rect 11093 2176 11095 2200
rect 11129 2200 11166 2210
rect 11129 2176 11131 2200
rect 11093 2166 11131 2176
rect 11165 2166 11166 2200
rect 10986 2142 11166 2166
rect 10986 2126 11023 2142
rect 10986 2092 10987 2126
rect 11021 2108 11023 2126
rect 11057 2126 11095 2142
rect 11057 2108 11059 2126
rect 11021 2092 11059 2108
rect 11093 2108 11095 2126
rect 11129 2126 11166 2142
rect 11129 2108 11131 2126
rect 11093 2092 11131 2108
rect 11165 2092 11166 2126
rect 10986 2074 11166 2092
rect 10986 2052 11023 2074
rect 10986 2018 10987 2052
rect 11021 2040 11023 2052
rect 11057 2052 11095 2074
rect 11057 2040 11059 2052
rect 11021 2018 11059 2040
rect 11093 2040 11095 2052
rect 11129 2052 11166 2074
rect 11129 2040 11131 2052
rect 11093 2018 11131 2040
rect 11165 2018 11166 2052
rect 10986 2006 11166 2018
rect 10986 1978 11023 2006
rect 10986 1944 10987 1978
rect 11021 1972 11023 1978
rect 11057 1978 11095 2006
rect 11057 1972 11059 1978
rect 11021 1944 11059 1972
rect 11093 1972 11095 1978
rect 11129 1978 11166 2006
rect 11129 1972 11131 1978
rect 11093 1944 11131 1972
rect 11165 1944 11166 1978
rect 10986 1938 11166 1944
rect 10986 1904 11023 1938
rect 11057 1904 11095 1938
rect 11129 1904 11166 1938
rect 10986 1870 10987 1904
rect 11021 1870 11059 1904
rect 11093 1870 11131 1904
rect 11165 1870 11166 1904
rect 10986 1836 11023 1870
rect 11057 1836 11095 1870
rect 11129 1836 11166 1870
rect 10986 1830 11166 1836
rect 10986 1796 10987 1830
rect 11021 1802 11059 1830
rect 11021 1796 11023 1802
rect 10986 1768 11023 1796
rect 11057 1796 11059 1802
rect 11093 1802 11131 1830
rect 11093 1796 11095 1802
rect 11057 1768 11095 1796
rect 11129 1796 11131 1802
rect 11165 1796 11166 1830
rect 11129 1768 11166 1796
rect 10986 1756 11166 1768
rect 10986 1722 10987 1756
rect 11021 1734 11059 1756
rect 11021 1722 11023 1734
rect 10986 1700 11023 1722
rect 11057 1722 11059 1734
rect 11093 1734 11131 1756
rect 11093 1722 11095 1734
rect 11057 1700 11095 1722
rect 11129 1722 11131 1734
rect 11165 1722 11166 1756
rect 11129 1700 11166 1722
rect 10986 1682 11166 1700
rect 10986 1648 10987 1682
rect 11021 1666 11059 1682
rect 11021 1648 11023 1666
rect 10986 1632 11023 1648
rect 11057 1648 11059 1666
rect 11093 1666 11131 1682
rect 11093 1648 11095 1666
rect 11057 1632 11095 1648
rect 11129 1648 11131 1666
rect 11165 1648 11166 1682
rect 11129 1632 11166 1648
rect 10986 1608 11166 1632
rect 10986 1574 10987 1608
rect 11021 1598 11059 1608
rect 11021 1574 11023 1598
rect 10986 1564 11023 1574
rect 11057 1574 11059 1598
rect 11093 1598 11131 1608
rect 11093 1574 11095 1598
rect 11057 1564 11095 1574
rect 11129 1574 11131 1598
rect 11165 1574 11166 1608
rect 11129 1564 11166 1574
rect 10986 1548 11166 1564
rect 11231 3104 11351 4200
rect 11793 4308 11913 4324
rect 11793 4274 11836 4308
rect 11870 4274 11913 4308
rect 11793 4234 11913 4274
rect 11793 4200 11836 4234
rect 11870 4200 11913 4234
rect 11231 3070 11274 3104
rect 11308 3070 11351 3104
rect 11231 3026 11351 3070
rect 11231 2992 11274 3026
rect 11308 2992 11351 3026
rect 11231 2948 11351 2992
rect 11231 2914 11274 2948
rect 11308 2914 11351 2948
rect 11231 2870 11351 2914
rect 11231 2836 11274 2870
rect 11308 2836 11351 2870
rect 11231 2792 11351 2836
rect 11231 2758 11274 2792
rect 11308 2758 11351 2792
rect 11231 2713 11351 2758
rect 11231 2679 11274 2713
rect 11308 2679 11351 2713
rect 11231 2634 11351 2679
rect 11231 2600 11274 2634
rect 11308 2600 11351 2634
rect 10801 1470 10844 1504
rect 10878 1470 10921 1504
rect 10801 1430 10921 1470
rect 10801 1396 10844 1430
rect 10878 1396 10921 1430
rect 10801 1250 10921 1396
rect 10801 1144 10808 1250
rect 10914 1144 10921 1250
rect 11231 1504 11351 2600
rect 11453 4092 11555 4118
rect 11589 4092 11691 4118
rect 11453 4082 11483 4092
rect 11661 4082 11691 4092
rect 11453 4014 11483 4048
rect 11661 4014 11691 4048
rect 11453 3946 11483 3980
rect 11661 3946 11691 3980
rect 11453 3878 11483 3912
rect 11661 3878 11691 3912
rect 11453 3810 11483 3844
rect 11661 3810 11691 3844
rect 11453 3742 11483 3776
rect 11661 3742 11691 3776
rect 11453 3674 11483 3708
rect 11661 3674 11691 3708
rect 11453 3606 11483 3640
rect 11661 3606 11691 3640
rect 11453 3538 11483 3572
rect 11661 3538 11691 3572
rect 11453 3470 11483 3504
rect 11661 3470 11691 3504
rect 11453 3402 11483 3436
rect 11661 3402 11691 3436
rect 11453 3334 11483 3368
rect 11661 3334 11691 3368
rect 11453 3266 11483 3300
rect 11661 3266 11691 3300
rect 11453 3198 11483 3232
rect 11661 3198 11691 3232
rect 11487 3164 11555 3194
rect 11589 3164 11657 3194
rect 11453 3148 11555 3164
rect 11589 3148 11691 3164
rect 11453 3108 11691 3148
rect 11453 3074 11483 3108
rect 11517 3074 11555 3108
rect 11589 3074 11627 3108
rect 11661 3074 11691 3108
rect 11453 3044 11691 3074
rect 11453 3028 11521 3044
rect 11453 2994 11483 3028
rect 11517 3010 11521 3028
rect 11555 3028 11589 3044
rect 11517 2994 11555 3010
rect 11623 3028 11691 3044
rect 11623 3010 11627 3028
rect 11589 2994 11627 3010
rect 11661 2994 11691 3028
rect 11453 2974 11691 2994
rect 11453 2948 11521 2974
rect 11453 2914 11483 2948
rect 11517 2940 11521 2948
rect 11555 2948 11589 2974
rect 11517 2914 11555 2940
rect 11623 2948 11691 2974
rect 11623 2940 11627 2948
rect 11589 2914 11627 2940
rect 11661 2914 11691 2948
rect 11453 2904 11691 2914
rect 11453 2870 11521 2904
rect 11555 2870 11589 2904
rect 11623 2870 11691 2904
rect 11453 2868 11691 2870
rect 11453 2834 11483 2868
rect 11517 2834 11555 2868
rect 11589 2834 11627 2868
rect 11661 2834 11691 2868
rect 11453 2800 11521 2834
rect 11555 2800 11589 2834
rect 11623 2800 11691 2834
rect 11453 2788 11691 2800
rect 11453 2754 11483 2788
rect 11517 2764 11555 2788
rect 11517 2754 11521 2764
rect 11453 2730 11521 2754
rect 11589 2764 11627 2788
rect 11555 2730 11589 2754
rect 11623 2754 11627 2764
rect 11661 2754 11691 2788
rect 11623 2730 11691 2754
rect 11453 2708 11691 2730
rect 11453 2674 11483 2708
rect 11517 2694 11555 2708
rect 11517 2674 11521 2694
rect 11453 2660 11521 2674
rect 11589 2694 11627 2708
rect 11555 2660 11589 2674
rect 11623 2674 11627 2694
rect 11661 2674 11691 2708
rect 11623 2660 11691 2674
rect 11453 2628 11691 2660
rect 11453 2594 11483 2628
rect 11517 2594 11555 2628
rect 11589 2594 11627 2628
rect 11661 2594 11691 2628
rect 11453 2556 11691 2594
rect 11453 2540 11555 2556
rect 11589 2540 11691 2556
rect 11487 2518 11555 2540
rect 11589 2518 11657 2540
rect 11453 2472 11483 2506
rect 11661 2472 11691 2506
rect 11453 2404 11483 2438
rect 11661 2404 11691 2438
rect 11453 2336 11483 2370
rect 11661 2336 11691 2370
rect 11453 2268 11483 2302
rect 11661 2268 11691 2302
rect 11453 2200 11483 2234
rect 11661 2200 11691 2234
rect 11453 2132 11483 2166
rect 11661 2132 11691 2166
rect 11453 2064 11483 2098
rect 11661 2064 11691 2098
rect 11453 1996 11483 2030
rect 11661 1996 11691 2030
rect 11453 1928 11483 1962
rect 11661 1928 11691 1962
rect 11453 1860 11483 1894
rect 11661 1860 11691 1894
rect 11453 1792 11483 1826
rect 11661 1792 11691 1826
rect 11453 1724 11483 1758
rect 11661 1724 11691 1758
rect 11453 1656 11483 1690
rect 11661 1656 11691 1690
rect 11453 1620 11483 1622
rect 11661 1620 11691 1622
rect 11453 1586 11555 1620
rect 11589 1586 11691 1620
rect 11453 1536 11691 1586
rect 11793 3104 11913 4200
rect 12223 4308 12343 4324
rect 12223 4274 12266 4308
rect 12300 4274 12343 4308
rect 12223 4234 12343 4274
rect 12223 4200 12266 4234
rect 12300 4200 12343 4234
rect 11793 3070 11836 3104
rect 11870 3070 11913 3104
rect 11793 3026 11913 3070
rect 11793 2992 11836 3026
rect 11870 2992 11913 3026
rect 11793 2948 11913 2992
rect 11793 2914 11836 2948
rect 11870 2914 11913 2948
rect 11793 2870 11913 2914
rect 11793 2836 11836 2870
rect 11870 2836 11913 2870
rect 11793 2792 11913 2836
rect 11793 2758 11836 2792
rect 11870 2758 11913 2792
rect 11793 2713 11913 2758
rect 11793 2679 11836 2713
rect 11870 2679 11913 2713
rect 11793 2634 11913 2679
rect 11793 2600 11836 2634
rect 11870 2600 11913 2634
rect 11231 1470 11274 1504
rect 11308 1470 11351 1504
rect 11231 1430 11351 1470
rect 11231 1396 11274 1430
rect 11308 1396 11351 1430
rect 11231 1250 11351 1396
rect 11231 1144 11238 1250
rect 11344 1144 11351 1250
rect 11793 1504 11913 2600
rect 11978 4064 11979 4098
rect 12013 4082 12051 4098
rect 12013 4064 12015 4082
rect 11978 4048 12015 4064
rect 12049 4064 12051 4082
rect 12085 4082 12123 4098
rect 12085 4064 12087 4082
rect 12049 4048 12087 4064
rect 12121 4064 12123 4082
rect 12157 4064 12158 4098
rect 12121 4048 12158 4064
rect 11978 4025 12158 4048
rect 11978 3991 11979 4025
rect 12013 4014 12051 4025
rect 12013 3991 12015 4014
rect 11978 3980 12015 3991
rect 12049 3991 12051 4014
rect 12085 4014 12123 4025
rect 12085 3991 12087 4014
rect 12049 3980 12087 3991
rect 12121 3991 12123 4014
rect 12157 3991 12158 4025
rect 12121 3980 12158 3991
rect 11978 3952 12158 3980
rect 11978 3918 11979 3952
rect 12013 3946 12051 3952
rect 12013 3918 12015 3946
rect 11978 3912 12015 3918
rect 12049 3918 12051 3946
rect 12085 3946 12123 3952
rect 12085 3918 12087 3946
rect 12049 3912 12087 3918
rect 12121 3918 12123 3946
rect 12157 3918 12158 3952
rect 12121 3912 12158 3918
rect 11978 3879 12158 3912
rect 11978 3845 11979 3879
rect 12013 3878 12051 3879
rect 12013 3845 12015 3878
rect 11978 3844 12015 3845
rect 12049 3845 12051 3878
rect 12085 3878 12123 3879
rect 12085 3845 12087 3878
rect 12049 3844 12087 3845
rect 12121 3845 12123 3878
rect 12157 3845 12158 3879
rect 12121 3844 12158 3845
rect 11978 3810 12158 3844
rect 11978 3806 12015 3810
rect 11978 3772 11979 3806
rect 12013 3776 12015 3806
rect 12049 3806 12087 3810
rect 12049 3776 12051 3806
rect 12013 3772 12051 3776
rect 12085 3776 12087 3806
rect 12121 3806 12158 3810
rect 12121 3776 12123 3806
rect 12085 3772 12123 3776
rect 12157 3772 12158 3806
rect 11978 3742 12158 3772
rect 11978 3733 12015 3742
rect 11978 3699 11979 3733
rect 12013 3708 12015 3733
rect 12049 3733 12087 3742
rect 12049 3708 12051 3733
rect 12013 3699 12051 3708
rect 12085 3708 12087 3733
rect 12121 3733 12158 3742
rect 12121 3708 12123 3733
rect 12085 3699 12123 3708
rect 12157 3699 12158 3733
rect 11978 3674 12158 3699
rect 11978 3660 12015 3674
rect 11978 3626 11979 3660
rect 12013 3640 12015 3660
rect 12049 3660 12087 3674
rect 12049 3640 12051 3660
rect 12013 3626 12051 3640
rect 12085 3640 12087 3660
rect 12121 3660 12158 3674
rect 12121 3640 12123 3660
rect 12085 3626 12123 3640
rect 12157 3626 12158 3660
rect 11978 3606 12158 3626
rect 11978 3587 12015 3606
rect 11978 3553 11979 3587
rect 12013 3572 12015 3587
rect 12049 3587 12087 3606
rect 12049 3572 12051 3587
rect 12013 3553 12051 3572
rect 12085 3572 12087 3587
rect 12121 3587 12158 3606
rect 12121 3572 12123 3587
rect 12085 3553 12123 3572
rect 12157 3553 12158 3587
rect 11978 3538 12158 3553
rect 11978 3514 12015 3538
rect 11978 3480 11979 3514
rect 12013 3504 12015 3514
rect 12049 3514 12087 3538
rect 12049 3504 12051 3514
rect 12013 3480 12051 3504
rect 12085 3504 12087 3514
rect 12121 3514 12158 3538
rect 12121 3504 12123 3514
rect 12085 3480 12123 3504
rect 12157 3480 12158 3514
rect 11978 3470 12158 3480
rect 11978 3441 12015 3470
rect 11978 3407 11979 3441
rect 12013 3436 12015 3441
rect 12049 3441 12087 3470
rect 12049 3436 12051 3441
rect 12013 3407 12051 3436
rect 12085 3436 12087 3441
rect 12121 3441 12158 3470
rect 12121 3436 12123 3441
rect 12085 3407 12123 3436
rect 12157 3407 12158 3441
rect 11978 3402 12158 3407
rect 11978 3368 12015 3402
rect 12049 3368 12087 3402
rect 12121 3368 12158 3402
rect 11978 3334 11979 3368
rect 12013 3334 12051 3368
rect 12085 3334 12123 3368
rect 12157 3334 12158 3368
rect 11978 3300 12015 3334
rect 12049 3300 12087 3334
rect 12121 3300 12158 3334
rect 11978 3295 12158 3300
rect 11978 3261 11979 3295
rect 12013 3266 12051 3295
rect 12013 3261 12015 3266
rect 11978 3232 12015 3261
rect 12049 3261 12051 3266
rect 12085 3266 12123 3295
rect 12085 3261 12087 3266
rect 12049 3232 12087 3261
rect 12121 3261 12123 3266
rect 12157 3261 12158 3295
rect 12121 3232 12158 3261
rect 11978 3222 12158 3232
rect 11978 3188 11979 3222
rect 12013 3198 12051 3222
rect 12013 3188 12015 3198
rect 11978 3164 12015 3188
rect 12049 3188 12051 3198
rect 12085 3198 12123 3222
rect 12085 3188 12087 3198
rect 12049 3164 12087 3188
rect 12121 3188 12123 3198
rect 12157 3188 12158 3222
rect 12121 3164 12158 3188
rect 11978 3149 12158 3164
rect 11978 3115 11979 3149
rect 12013 3115 12051 3149
rect 12085 3115 12123 3149
rect 12157 3115 12158 3149
rect 11978 3076 12158 3115
rect 11978 3042 11979 3076
rect 12013 3042 12051 3076
rect 12085 3042 12123 3076
rect 12157 3042 12158 3076
rect 11978 3003 12158 3042
rect 11978 2969 11979 3003
rect 12013 2969 12051 3003
rect 12085 2969 12123 3003
rect 12157 2969 12158 3003
rect 11978 2930 12158 2969
rect 11978 2896 11979 2930
rect 12013 2896 12051 2930
rect 12085 2896 12123 2930
rect 12157 2896 12158 2930
rect 11978 2857 12158 2896
rect 11978 2823 11979 2857
rect 12013 2823 12051 2857
rect 12085 2823 12123 2857
rect 12157 2823 12158 2857
rect 11978 2784 12158 2823
rect 11978 2750 11979 2784
rect 12013 2750 12051 2784
rect 12085 2750 12123 2784
rect 12157 2750 12158 2784
rect 11978 2711 12158 2750
rect 11978 2677 11979 2711
rect 12013 2677 12051 2711
rect 12085 2677 12123 2711
rect 12157 2677 12158 2711
rect 11978 2638 12158 2677
rect 11978 2604 11979 2638
rect 12013 2604 12051 2638
rect 12085 2604 12123 2638
rect 12157 2604 12158 2638
rect 11978 2565 12158 2604
rect 11978 2531 11979 2565
rect 12013 2531 12051 2565
rect 12085 2531 12123 2565
rect 12157 2531 12158 2565
rect 11978 2492 12158 2531
rect 11978 2458 11979 2492
rect 12013 2482 12051 2492
rect 12013 2458 12015 2482
rect 11978 2448 12015 2458
rect 12049 2458 12051 2482
rect 12085 2482 12123 2492
rect 12085 2458 12087 2482
rect 12049 2448 12087 2458
rect 12121 2458 12123 2482
rect 12157 2458 12158 2492
rect 12121 2448 12158 2458
rect 11978 2419 12158 2448
rect 11978 2385 11979 2419
rect 12013 2414 12051 2419
rect 12013 2385 12015 2414
rect 11978 2380 12015 2385
rect 12049 2385 12051 2414
rect 12085 2414 12123 2419
rect 12085 2385 12087 2414
rect 12049 2380 12087 2385
rect 12121 2385 12123 2414
rect 12157 2385 12158 2419
rect 12121 2380 12158 2385
rect 11978 2346 12158 2380
rect 11978 2312 11979 2346
rect 12013 2312 12015 2346
rect 12049 2312 12051 2346
rect 12085 2312 12087 2346
rect 12121 2312 12123 2346
rect 12157 2312 12158 2346
rect 11978 2278 12158 2312
rect 11978 2273 12015 2278
rect 11978 2239 11979 2273
rect 12013 2244 12015 2273
rect 12049 2273 12087 2278
rect 12049 2244 12051 2273
rect 12013 2239 12051 2244
rect 12085 2244 12087 2273
rect 12121 2273 12158 2278
rect 12121 2244 12123 2273
rect 12085 2239 12123 2244
rect 12157 2239 12158 2273
rect 11978 2210 12158 2239
rect 11978 2200 12015 2210
rect 11978 2166 11979 2200
rect 12013 2176 12015 2200
rect 12049 2200 12087 2210
rect 12049 2176 12051 2200
rect 12013 2166 12051 2176
rect 12085 2176 12087 2200
rect 12121 2200 12158 2210
rect 12121 2176 12123 2200
rect 12085 2166 12123 2176
rect 12157 2166 12158 2200
rect 11978 2142 12158 2166
rect 11978 2126 12015 2142
rect 11978 2092 11979 2126
rect 12013 2108 12015 2126
rect 12049 2126 12087 2142
rect 12049 2108 12051 2126
rect 12013 2092 12051 2108
rect 12085 2108 12087 2126
rect 12121 2126 12158 2142
rect 12121 2108 12123 2126
rect 12085 2092 12123 2108
rect 12157 2092 12158 2126
rect 11978 2074 12158 2092
rect 11978 2052 12015 2074
rect 11978 2018 11979 2052
rect 12013 2040 12015 2052
rect 12049 2052 12087 2074
rect 12049 2040 12051 2052
rect 12013 2018 12051 2040
rect 12085 2040 12087 2052
rect 12121 2052 12158 2074
rect 12121 2040 12123 2052
rect 12085 2018 12123 2040
rect 12157 2018 12158 2052
rect 11978 2006 12158 2018
rect 11978 1978 12015 2006
rect 11978 1944 11979 1978
rect 12013 1972 12015 1978
rect 12049 1978 12087 2006
rect 12049 1972 12051 1978
rect 12013 1944 12051 1972
rect 12085 1972 12087 1978
rect 12121 1978 12158 2006
rect 12121 1972 12123 1978
rect 12085 1944 12123 1972
rect 12157 1944 12158 1978
rect 11978 1938 12158 1944
rect 11978 1904 12015 1938
rect 12049 1904 12087 1938
rect 12121 1904 12158 1938
rect 11978 1870 11979 1904
rect 12013 1870 12051 1904
rect 12085 1870 12123 1904
rect 12157 1870 12158 1904
rect 11978 1836 12015 1870
rect 12049 1836 12087 1870
rect 12121 1836 12158 1870
rect 11978 1830 12158 1836
rect 11978 1796 11979 1830
rect 12013 1802 12051 1830
rect 12013 1796 12015 1802
rect 11978 1768 12015 1796
rect 12049 1796 12051 1802
rect 12085 1802 12123 1830
rect 12085 1796 12087 1802
rect 12049 1768 12087 1796
rect 12121 1796 12123 1802
rect 12157 1796 12158 1830
rect 12121 1768 12158 1796
rect 11978 1756 12158 1768
rect 11978 1722 11979 1756
rect 12013 1734 12051 1756
rect 12013 1722 12015 1734
rect 11978 1700 12015 1722
rect 12049 1722 12051 1734
rect 12085 1734 12123 1756
rect 12085 1722 12087 1734
rect 12049 1700 12087 1722
rect 12121 1722 12123 1734
rect 12157 1722 12158 1756
rect 12121 1700 12158 1722
rect 11978 1682 12158 1700
rect 11978 1648 11979 1682
rect 12013 1666 12051 1682
rect 12013 1648 12015 1666
rect 11978 1632 12015 1648
rect 12049 1648 12051 1666
rect 12085 1666 12123 1682
rect 12085 1648 12087 1666
rect 12049 1632 12087 1648
rect 12121 1648 12123 1666
rect 12157 1648 12158 1682
rect 12121 1632 12158 1648
rect 11978 1608 12158 1632
rect 11978 1574 11979 1608
rect 12013 1598 12051 1608
rect 12013 1574 12015 1598
rect 11978 1564 12015 1574
rect 12049 1574 12051 1598
rect 12085 1598 12123 1608
rect 12085 1574 12087 1598
rect 12049 1564 12087 1574
rect 12121 1574 12123 1598
rect 12157 1574 12158 1608
rect 12121 1564 12158 1574
rect 11978 1548 12158 1564
rect 12223 3104 12343 4200
rect 12785 4308 12905 4324
rect 12785 4274 12828 4308
rect 12862 4274 12905 4308
rect 12785 4234 12905 4274
rect 12785 4200 12828 4234
rect 12862 4200 12905 4234
rect 12223 3070 12266 3104
rect 12300 3070 12343 3104
rect 12223 3026 12343 3070
rect 12223 2992 12266 3026
rect 12300 2992 12343 3026
rect 12223 2948 12343 2992
rect 12223 2914 12266 2948
rect 12300 2914 12343 2948
rect 12223 2870 12343 2914
rect 12223 2836 12266 2870
rect 12300 2836 12343 2870
rect 12223 2792 12343 2836
rect 12223 2758 12266 2792
rect 12300 2758 12343 2792
rect 12223 2713 12343 2758
rect 12223 2679 12266 2713
rect 12300 2679 12343 2713
rect 12223 2634 12343 2679
rect 12223 2600 12266 2634
rect 12300 2600 12343 2634
rect 11793 1470 11836 1504
rect 11870 1470 11913 1504
rect 11793 1430 11913 1470
rect 11793 1396 11836 1430
rect 11870 1396 11913 1430
rect 11793 1250 11913 1396
rect 11793 1144 11800 1250
rect 11906 1144 11913 1250
rect 12223 1504 12343 2600
rect 12445 4092 12547 4118
rect 12581 4092 12683 4118
rect 12445 4082 12475 4092
rect 12653 4082 12683 4092
rect 12445 4014 12475 4048
rect 12653 4014 12683 4048
rect 12445 3946 12475 3980
rect 12653 3946 12683 3980
rect 12445 3878 12475 3912
rect 12653 3878 12683 3912
rect 12445 3810 12475 3844
rect 12653 3810 12683 3844
rect 12445 3742 12475 3776
rect 12653 3742 12683 3776
rect 12445 3674 12475 3708
rect 12653 3674 12683 3708
rect 12445 3606 12475 3640
rect 12653 3606 12683 3640
rect 12445 3538 12475 3572
rect 12653 3538 12683 3572
rect 12445 3470 12475 3504
rect 12653 3470 12683 3504
rect 12445 3402 12475 3436
rect 12653 3402 12683 3436
rect 12445 3334 12475 3368
rect 12653 3334 12683 3368
rect 12445 3266 12475 3300
rect 12653 3266 12683 3300
rect 12445 3198 12475 3232
rect 12653 3198 12683 3232
rect 12479 3164 12547 3194
rect 12581 3164 12649 3194
rect 12445 3148 12547 3164
rect 12581 3148 12683 3164
rect 12445 3108 12683 3148
rect 12445 3074 12475 3108
rect 12509 3074 12547 3108
rect 12581 3074 12619 3108
rect 12653 3074 12683 3108
rect 12445 3044 12683 3074
rect 12445 3028 12513 3044
rect 12445 2994 12475 3028
rect 12509 3010 12513 3028
rect 12547 3028 12581 3044
rect 12509 2994 12547 3010
rect 12615 3028 12683 3044
rect 12615 3010 12619 3028
rect 12581 2994 12619 3010
rect 12653 2994 12683 3028
rect 12445 2974 12683 2994
rect 12445 2948 12513 2974
rect 12445 2914 12475 2948
rect 12509 2940 12513 2948
rect 12547 2948 12581 2974
rect 12509 2914 12547 2940
rect 12615 2948 12683 2974
rect 12615 2940 12619 2948
rect 12581 2914 12619 2940
rect 12653 2914 12683 2948
rect 12445 2904 12683 2914
rect 12445 2870 12513 2904
rect 12547 2870 12581 2904
rect 12615 2870 12683 2904
rect 12445 2868 12683 2870
rect 12445 2834 12475 2868
rect 12509 2834 12547 2868
rect 12581 2834 12619 2868
rect 12653 2834 12683 2868
rect 12445 2800 12513 2834
rect 12547 2800 12581 2834
rect 12615 2800 12683 2834
rect 12445 2788 12683 2800
rect 12445 2754 12475 2788
rect 12509 2764 12547 2788
rect 12509 2754 12513 2764
rect 12445 2730 12513 2754
rect 12581 2764 12619 2788
rect 12547 2730 12581 2754
rect 12615 2754 12619 2764
rect 12653 2754 12683 2788
rect 12615 2730 12683 2754
rect 12445 2708 12683 2730
rect 12445 2674 12475 2708
rect 12509 2694 12547 2708
rect 12509 2674 12513 2694
rect 12445 2660 12513 2674
rect 12581 2694 12619 2708
rect 12547 2660 12581 2674
rect 12615 2674 12619 2694
rect 12653 2674 12683 2708
rect 12615 2660 12683 2674
rect 12445 2628 12683 2660
rect 12445 2594 12475 2628
rect 12509 2594 12547 2628
rect 12581 2594 12619 2628
rect 12653 2594 12683 2628
rect 12445 2556 12683 2594
rect 12445 2540 12547 2556
rect 12581 2540 12683 2556
rect 12479 2518 12547 2540
rect 12581 2518 12649 2540
rect 12445 2472 12475 2506
rect 12653 2472 12683 2506
rect 12445 2404 12475 2438
rect 12653 2404 12683 2438
rect 12445 2336 12475 2370
rect 12653 2336 12683 2370
rect 12445 2268 12475 2302
rect 12653 2268 12683 2302
rect 12445 2200 12475 2234
rect 12653 2200 12683 2234
rect 12445 2132 12475 2166
rect 12653 2132 12683 2166
rect 12445 2064 12475 2098
rect 12653 2064 12683 2098
rect 12445 1996 12475 2030
rect 12653 1996 12683 2030
rect 12445 1928 12475 1962
rect 12653 1928 12683 1962
rect 12445 1860 12475 1894
rect 12653 1860 12683 1894
rect 12445 1792 12475 1826
rect 12653 1792 12683 1826
rect 12445 1724 12475 1758
rect 12653 1724 12683 1758
rect 12445 1656 12475 1690
rect 12653 1656 12683 1690
rect 12445 1620 12475 1622
rect 12653 1620 12683 1622
rect 12445 1586 12547 1620
rect 12581 1586 12683 1620
rect 12445 1536 12683 1586
rect 12785 3104 12905 4200
rect 13215 4308 13335 4324
rect 13215 4274 13258 4308
rect 13292 4274 13335 4308
rect 13215 4234 13335 4274
rect 13215 4200 13258 4234
rect 13292 4200 13335 4234
rect 12785 3070 12828 3104
rect 12862 3070 12905 3104
rect 12785 3026 12905 3070
rect 12785 2992 12828 3026
rect 12862 2992 12905 3026
rect 12785 2948 12905 2992
rect 12785 2914 12828 2948
rect 12862 2914 12905 2948
rect 12785 2870 12905 2914
rect 12785 2836 12828 2870
rect 12862 2836 12905 2870
rect 12785 2792 12905 2836
rect 12785 2758 12828 2792
rect 12862 2758 12905 2792
rect 12785 2713 12905 2758
rect 12785 2679 12828 2713
rect 12862 2679 12905 2713
rect 12785 2634 12905 2679
rect 12785 2600 12828 2634
rect 12862 2600 12905 2634
rect 12223 1470 12266 1504
rect 12300 1470 12343 1504
rect 12223 1430 12343 1470
rect 12223 1396 12266 1430
rect 12300 1396 12343 1430
rect 12223 1250 12343 1396
rect 12223 1144 12230 1250
rect 12336 1144 12343 1250
rect 12785 1504 12905 2600
rect 12970 4064 12971 4098
rect 13005 4082 13043 4098
rect 13005 4064 13007 4082
rect 12970 4048 13007 4064
rect 13041 4064 13043 4082
rect 13077 4082 13115 4098
rect 13077 4064 13079 4082
rect 13041 4048 13079 4064
rect 13113 4064 13115 4082
rect 13149 4064 13150 4098
rect 13113 4048 13150 4064
rect 12970 4025 13150 4048
rect 12970 3991 12971 4025
rect 13005 4014 13043 4025
rect 13005 3991 13007 4014
rect 12970 3980 13007 3991
rect 13041 3991 13043 4014
rect 13077 4014 13115 4025
rect 13077 3991 13079 4014
rect 13041 3980 13079 3991
rect 13113 3991 13115 4014
rect 13149 3991 13150 4025
rect 13113 3980 13150 3991
rect 12970 3952 13150 3980
rect 12970 3918 12971 3952
rect 13005 3946 13043 3952
rect 13005 3918 13007 3946
rect 12970 3912 13007 3918
rect 13041 3918 13043 3946
rect 13077 3946 13115 3952
rect 13077 3918 13079 3946
rect 13041 3912 13079 3918
rect 13113 3918 13115 3946
rect 13149 3918 13150 3952
rect 13113 3912 13150 3918
rect 12970 3879 13150 3912
rect 12970 3845 12971 3879
rect 13005 3878 13043 3879
rect 13005 3845 13007 3878
rect 12970 3844 13007 3845
rect 13041 3845 13043 3878
rect 13077 3878 13115 3879
rect 13077 3845 13079 3878
rect 13041 3844 13079 3845
rect 13113 3845 13115 3878
rect 13149 3845 13150 3879
rect 13113 3844 13150 3845
rect 12970 3810 13150 3844
rect 12970 3806 13007 3810
rect 12970 3772 12971 3806
rect 13005 3776 13007 3806
rect 13041 3806 13079 3810
rect 13041 3776 13043 3806
rect 13005 3772 13043 3776
rect 13077 3776 13079 3806
rect 13113 3806 13150 3810
rect 13113 3776 13115 3806
rect 13077 3772 13115 3776
rect 13149 3772 13150 3806
rect 12970 3742 13150 3772
rect 12970 3733 13007 3742
rect 12970 3699 12971 3733
rect 13005 3708 13007 3733
rect 13041 3733 13079 3742
rect 13041 3708 13043 3733
rect 13005 3699 13043 3708
rect 13077 3708 13079 3733
rect 13113 3733 13150 3742
rect 13113 3708 13115 3733
rect 13077 3699 13115 3708
rect 13149 3699 13150 3733
rect 12970 3674 13150 3699
rect 12970 3660 13007 3674
rect 12970 3626 12971 3660
rect 13005 3640 13007 3660
rect 13041 3660 13079 3674
rect 13041 3640 13043 3660
rect 13005 3626 13043 3640
rect 13077 3640 13079 3660
rect 13113 3660 13150 3674
rect 13113 3640 13115 3660
rect 13077 3626 13115 3640
rect 13149 3626 13150 3660
rect 12970 3606 13150 3626
rect 12970 3587 13007 3606
rect 12970 3553 12971 3587
rect 13005 3572 13007 3587
rect 13041 3587 13079 3606
rect 13041 3572 13043 3587
rect 13005 3553 13043 3572
rect 13077 3572 13079 3587
rect 13113 3587 13150 3606
rect 13113 3572 13115 3587
rect 13077 3553 13115 3572
rect 13149 3553 13150 3587
rect 12970 3538 13150 3553
rect 12970 3514 13007 3538
rect 12970 3480 12971 3514
rect 13005 3504 13007 3514
rect 13041 3514 13079 3538
rect 13041 3504 13043 3514
rect 13005 3480 13043 3504
rect 13077 3504 13079 3514
rect 13113 3514 13150 3538
rect 13113 3504 13115 3514
rect 13077 3480 13115 3504
rect 13149 3480 13150 3514
rect 12970 3470 13150 3480
rect 12970 3441 13007 3470
rect 12970 3407 12971 3441
rect 13005 3436 13007 3441
rect 13041 3441 13079 3470
rect 13041 3436 13043 3441
rect 13005 3407 13043 3436
rect 13077 3436 13079 3441
rect 13113 3441 13150 3470
rect 13113 3436 13115 3441
rect 13077 3407 13115 3436
rect 13149 3407 13150 3441
rect 12970 3402 13150 3407
rect 12970 3368 13007 3402
rect 13041 3368 13079 3402
rect 13113 3368 13150 3402
rect 12970 3334 12971 3368
rect 13005 3334 13043 3368
rect 13077 3334 13115 3368
rect 13149 3334 13150 3368
rect 12970 3300 13007 3334
rect 13041 3300 13079 3334
rect 13113 3300 13150 3334
rect 12970 3295 13150 3300
rect 12970 3261 12971 3295
rect 13005 3266 13043 3295
rect 13005 3261 13007 3266
rect 12970 3232 13007 3261
rect 13041 3261 13043 3266
rect 13077 3266 13115 3295
rect 13077 3261 13079 3266
rect 13041 3232 13079 3261
rect 13113 3261 13115 3266
rect 13149 3261 13150 3295
rect 13113 3232 13150 3261
rect 12970 3222 13150 3232
rect 12970 3188 12971 3222
rect 13005 3198 13043 3222
rect 13005 3188 13007 3198
rect 12970 3164 13007 3188
rect 13041 3188 13043 3198
rect 13077 3198 13115 3222
rect 13077 3188 13079 3198
rect 13041 3164 13079 3188
rect 13113 3188 13115 3198
rect 13149 3188 13150 3222
rect 13113 3164 13150 3188
rect 12970 3149 13150 3164
rect 12970 3115 12971 3149
rect 13005 3115 13043 3149
rect 13077 3115 13115 3149
rect 13149 3115 13150 3149
rect 12970 3076 13150 3115
rect 12970 3042 12971 3076
rect 13005 3042 13043 3076
rect 13077 3042 13115 3076
rect 13149 3042 13150 3076
rect 12970 3003 13150 3042
rect 12970 2969 12971 3003
rect 13005 2969 13043 3003
rect 13077 2969 13115 3003
rect 13149 2969 13150 3003
rect 12970 2930 13150 2969
rect 12970 2896 12971 2930
rect 13005 2896 13043 2930
rect 13077 2896 13115 2930
rect 13149 2896 13150 2930
rect 12970 2857 13150 2896
rect 12970 2823 12971 2857
rect 13005 2823 13043 2857
rect 13077 2823 13115 2857
rect 13149 2823 13150 2857
rect 12970 2784 13150 2823
rect 12970 2750 12971 2784
rect 13005 2750 13043 2784
rect 13077 2750 13115 2784
rect 13149 2750 13150 2784
rect 12970 2711 13150 2750
rect 12970 2677 12971 2711
rect 13005 2677 13043 2711
rect 13077 2677 13115 2711
rect 13149 2677 13150 2711
rect 12970 2638 13150 2677
rect 12970 2604 12971 2638
rect 13005 2604 13043 2638
rect 13077 2604 13115 2638
rect 13149 2604 13150 2638
rect 12970 2565 13150 2604
rect 12970 2531 12971 2565
rect 13005 2531 13043 2565
rect 13077 2531 13115 2565
rect 13149 2531 13150 2565
rect 12970 2492 13150 2531
rect 12970 2458 12971 2492
rect 13005 2482 13043 2492
rect 13005 2458 13007 2482
rect 12970 2448 13007 2458
rect 13041 2458 13043 2482
rect 13077 2482 13115 2492
rect 13077 2458 13079 2482
rect 13041 2448 13079 2458
rect 13113 2458 13115 2482
rect 13149 2458 13150 2492
rect 13113 2448 13150 2458
rect 12970 2419 13150 2448
rect 12970 2385 12971 2419
rect 13005 2414 13043 2419
rect 13005 2385 13007 2414
rect 12970 2380 13007 2385
rect 13041 2385 13043 2414
rect 13077 2414 13115 2419
rect 13077 2385 13079 2414
rect 13041 2380 13079 2385
rect 13113 2385 13115 2414
rect 13149 2385 13150 2419
rect 13113 2380 13150 2385
rect 12970 2346 13150 2380
rect 12970 2312 12971 2346
rect 13005 2312 13007 2346
rect 13041 2312 13043 2346
rect 13077 2312 13079 2346
rect 13113 2312 13115 2346
rect 13149 2312 13150 2346
rect 12970 2278 13150 2312
rect 12970 2273 13007 2278
rect 12970 2239 12971 2273
rect 13005 2244 13007 2273
rect 13041 2273 13079 2278
rect 13041 2244 13043 2273
rect 13005 2239 13043 2244
rect 13077 2244 13079 2273
rect 13113 2273 13150 2278
rect 13113 2244 13115 2273
rect 13077 2239 13115 2244
rect 13149 2239 13150 2273
rect 12970 2210 13150 2239
rect 12970 2200 13007 2210
rect 12970 2166 12971 2200
rect 13005 2176 13007 2200
rect 13041 2200 13079 2210
rect 13041 2176 13043 2200
rect 13005 2166 13043 2176
rect 13077 2176 13079 2200
rect 13113 2200 13150 2210
rect 13113 2176 13115 2200
rect 13077 2166 13115 2176
rect 13149 2166 13150 2200
rect 12970 2142 13150 2166
rect 12970 2126 13007 2142
rect 12970 2092 12971 2126
rect 13005 2108 13007 2126
rect 13041 2126 13079 2142
rect 13041 2108 13043 2126
rect 13005 2092 13043 2108
rect 13077 2108 13079 2126
rect 13113 2126 13150 2142
rect 13113 2108 13115 2126
rect 13077 2092 13115 2108
rect 13149 2092 13150 2126
rect 12970 2074 13150 2092
rect 12970 2052 13007 2074
rect 12970 2018 12971 2052
rect 13005 2040 13007 2052
rect 13041 2052 13079 2074
rect 13041 2040 13043 2052
rect 13005 2018 13043 2040
rect 13077 2040 13079 2052
rect 13113 2052 13150 2074
rect 13113 2040 13115 2052
rect 13077 2018 13115 2040
rect 13149 2018 13150 2052
rect 12970 2006 13150 2018
rect 12970 1978 13007 2006
rect 12970 1944 12971 1978
rect 13005 1972 13007 1978
rect 13041 1978 13079 2006
rect 13041 1972 13043 1978
rect 13005 1944 13043 1972
rect 13077 1972 13079 1978
rect 13113 1978 13150 2006
rect 13113 1972 13115 1978
rect 13077 1944 13115 1972
rect 13149 1944 13150 1978
rect 12970 1938 13150 1944
rect 12970 1904 13007 1938
rect 13041 1904 13079 1938
rect 13113 1904 13150 1938
rect 12970 1870 12971 1904
rect 13005 1870 13043 1904
rect 13077 1870 13115 1904
rect 13149 1870 13150 1904
rect 12970 1836 13007 1870
rect 13041 1836 13079 1870
rect 13113 1836 13150 1870
rect 12970 1830 13150 1836
rect 12970 1796 12971 1830
rect 13005 1802 13043 1830
rect 13005 1796 13007 1802
rect 12970 1768 13007 1796
rect 13041 1796 13043 1802
rect 13077 1802 13115 1830
rect 13077 1796 13079 1802
rect 13041 1768 13079 1796
rect 13113 1796 13115 1802
rect 13149 1796 13150 1830
rect 13113 1768 13150 1796
rect 12970 1756 13150 1768
rect 12970 1722 12971 1756
rect 13005 1734 13043 1756
rect 13005 1722 13007 1734
rect 12970 1700 13007 1722
rect 13041 1722 13043 1734
rect 13077 1734 13115 1756
rect 13077 1722 13079 1734
rect 13041 1700 13079 1722
rect 13113 1722 13115 1734
rect 13149 1722 13150 1756
rect 13113 1700 13150 1722
rect 12970 1682 13150 1700
rect 12970 1648 12971 1682
rect 13005 1666 13043 1682
rect 13005 1648 13007 1666
rect 12970 1632 13007 1648
rect 13041 1648 13043 1666
rect 13077 1666 13115 1682
rect 13077 1648 13079 1666
rect 13041 1632 13079 1648
rect 13113 1648 13115 1666
rect 13149 1648 13150 1682
rect 13113 1632 13150 1648
rect 12970 1608 13150 1632
rect 12970 1574 12971 1608
rect 13005 1598 13043 1608
rect 13005 1574 13007 1598
rect 12970 1564 13007 1574
rect 13041 1574 13043 1598
rect 13077 1598 13115 1608
rect 13077 1574 13079 1598
rect 13041 1564 13079 1574
rect 13113 1574 13115 1598
rect 13149 1574 13150 1608
rect 13113 1564 13150 1574
rect 12970 1548 13150 1564
rect 13215 3104 13335 4200
rect 13777 4308 13897 4324
rect 13777 4274 13820 4308
rect 13854 4274 13897 4308
rect 13777 4234 13897 4274
rect 13777 4200 13820 4234
rect 13854 4200 13897 4234
rect 13215 3070 13258 3104
rect 13292 3070 13335 3104
rect 13215 3026 13335 3070
rect 13215 2992 13258 3026
rect 13292 2992 13335 3026
rect 13215 2948 13335 2992
rect 13215 2914 13258 2948
rect 13292 2914 13335 2948
rect 13215 2870 13335 2914
rect 13215 2836 13258 2870
rect 13292 2836 13335 2870
rect 13215 2792 13335 2836
rect 13215 2758 13258 2792
rect 13292 2758 13335 2792
rect 13215 2713 13335 2758
rect 13215 2679 13258 2713
rect 13292 2679 13335 2713
rect 13215 2634 13335 2679
rect 13215 2600 13258 2634
rect 13292 2600 13335 2634
rect 12785 1470 12828 1504
rect 12862 1470 12905 1504
rect 12785 1430 12905 1470
rect 12785 1396 12828 1430
rect 12862 1396 12905 1430
rect 12785 1250 12905 1396
rect 12785 1144 12792 1250
rect 12898 1144 12905 1250
rect 13215 1504 13335 2600
rect 13437 4092 13539 4118
rect 13573 4092 13675 4118
rect 13437 4082 13467 4092
rect 13645 4082 13675 4092
rect 13437 4014 13467 4048
rect 13645 4014 13675 4048
rect 13437 3946 13467 3980
rect 13645 3946 13675 3980
rect 13437 3878 13467 3912
rect 13645 3878 13675 3912
rect 13437 3810 13467 3844
rect 13645 3810 13675 3844
rect 13437 3742 13467 3776
rect 13645 3742 13675 3776
rect 13437 3674 13467 3708
rect 13645 3674 13675 3708
rect 13437 3606 13467 3640
rect 13645 3606 13675 3640
rect 13437 3538 13467 3572
rect 13645 3538 13675 3572
rect 13437 3470 13467 3504
rect 13645 3470 13675 3504
rect 13437 3402 13467 3436
rect 13645 3402 13675 3436
rect 13437 3334 13467 3368
rect 13645 3334 13675 3368
rect 13437 3266 13467 3300
rect 13645 3266 13675 3300
rect 13437 3198 13467 3232
rect 13645 3198 13675 3232
rect 13471 3164 13539 3194
rect 13573 3164 13641 3194
rect 13437 3148 13539 3164
rect 13573 3148 13675 3164
rect 13437 3108 13675 3148
rect 13437 3074 13467 3108
rect 13501 3074 13539 3108
rect 13573 3074 13611 3108
rect 13645 3074 13675 3108
rect 13437 3044 13675 3074
rect 13437 3028 13505 3044
rect 13437 2994 13467 3028
rect 13501 3010 13505 3028
rect 13539 3028 13573 3044
rect 13501 2994 13539 3010
rect 13607 3028 13675 3044
rect 13607 3010 13611 3028
rect 13573 2994 13611 3010
rect 13645 2994 13675 3028
rect 13437 2974 13675 2994
rect 13437 2948 13505 2974
rect 13437 2914 13467 2948
rect 13501 2940 13505 2948
rect 13539 2948 13573 2974
rect 13501 2914 13539 2940
rect 13607 2948 13675 2974
rect 13607 2940 13611 2948
rect 13573 2914 13611 2940
rect 13645 2914 13675 2948
rect 13437 2904 13675 2914
rect 13437 2870 13505 2904
rect 13539 2870 13573 2904
rect 13607 2870 13675 2904
rect 13437 2868 13675 2870
rect 13437 2834 13467 2868
rect 13501 2834 13539 2868
rect 13573 2834 13611 2868
rect 13645 2834 13675 2868
rect 13437 2800 13505 2834
rect 13539 2800 13573 2834
rect 13607 2800 13675 2834
rect 13437 2788 13675 2800
rect 13437 2754 13467 2788
rect 13501 2764 13539 2788
rect 13501 2754 13505 2764
rect 13437 2730 13505 2754
rect 13573 2764 13611 2788
rect 13539 2730 13573 2754
rect 13607 2754 13611 2764
rect 13645 2754 13675 2788
rect 13607 2730 13675 2754
rect 13437 2708 13675 2730
rect 13437 2674 13467 2708
rect 13501 2694 13539 2708
rect 13501 2674 13505 2694
rect 13437 2660 13505 2674
rect 13573 2694 13611 2708
rect 13539 2660 13573 2674
rect 13607 2674 13611 2694
rect 13645 2674 13675 2708
rect 13607 2660 13675 2674
rect 13437 2628 13675 2660
rect 13437 2594 13467 2628
rect 13501 2594 13539 2628
rect 13573 2594 13611 2628
rect 13645 2594 13675 2628
rect 13437 2556 13675 2594
rect 13437 2540 13539 2556
rect 13573 2540 13675 2556
rect 13471 2518 13539 2540
rect 13573 2518 13641 2540
rect 13437 2472 13467 2506
rect 13645 2472 13675 2506
rect 13437 2404 13467 2438
rect 13645 2404 13675 2438
rect 13437 2336 13467 2370
rect 13645 2336 13675 2370
rect 13437 2268 13467 2302
rect 13645 2268 13675 2302
rect 13437 2200 13467 2234
rect 13645 2200 13675 2234
rect 13437 2132 13467 2166
rect 13645 2132 13675 2166
rect 13437 2064 13467 2098
rect 13645 2064 13675 2098
rect 13437 1996 13467 2030
rect 13645 1996 13675 2030
rect 13437 1928 13467 1962
rect 13645 1928 13675 1962
rect 13437 1860 13467 1894
rect 13645 1860 13675 1894
rect 13437 1792 13467 1826
rect 13645 1792 13675 1826
rect 13437 1724 13467 1758
rect 13645 1724 13675 1758
rect 13437 1656 13467 1690
rect 13645 1656 13675 1690
rect 13437 1620 13467 1622
rect 13645 1620 13675 1622
rect 13437 1586 13539 1620
rect 13573 1586 13675 1620
rect 13437 1536 13675 1586
rect 13777 3104 13897 4200
rect 14135 4308 14255 4324
rect 14135 4274 14178 4308
rect 14212 4274 14255 4308
rect 14135 4234 14255 4274
rect 14135 4200 14178 4234
rect 14212 4200 14255 4234
rect 13777 3070 13820 3104
rect 13854 3070 13897 3104
rect 13777 3026 13897 3070
rect 13777 2992 13820 3026
rect 13854 2992 13897 3026
rect 13777 2948 13897 2992
rect 13777 2914 13820 2948
rect 13854 2914 13897 2948
rect 13777 2870 13897 2914
rect 13777 2836 13820 2870
rect 13854 2836 13897 2870
rect 13777 2792 13897 2836
rect 13777 2758 13820 2792
rect 13854 2758 13897 2792
rect 13777 2713 13897 2758
rect 13777 2679 13820 2713
rect 13854 2679 13897 2713
rect 13777 2634 13897 2679
rect 13777 2600 13820 2634
rect 13854 2600 13897 2634
rect 13215 1470 13258 1504
rect 13292 1470 13335 1504
rect 13215 1430 13335 1470
rect 13215 1396 13258 1430
rect 13292 1396 13335 1430
rect 13215 1250 13335 1396
rect 13215 1144 13222 1250
rect 13328 1144 13335 1250
rect 13777 1504 13897 2600
rect 13999 4025 14033 4048
rect 13999 3952 14033 3980
rect 13999 3879 14033 3912
rect 13999 3810 14033 3844
rect 13999 3742 14033 3772
rect 13999 3674 14033 3699
rect 13999 3606 14033 3626
rect 13999 3538 14033 3553
rect 13999 3470 14033 3480
rect 13999 3402 14033 3407
rect 13999 3295 14033 3300
rect 13999 3222 14033 3232
rect 13999 3149 14033 3164
rect 13999 3076 14033 3115
rect 13999 3003 14033 3042
rect 13999 2930 14033 2969
rect 13999 2857 14033 2896
rect 13999 2784 14033 2823
rect 13999 2711 14033 2750
rect 13999 2638 14033 2677
rect 13999 2565 14033 2604
rect 13999 2492 14033 2531
rect 13999 2419 14033 2448
rect 13999 2346 14033 2380
rect 13999 2278 14033 2312
rect 13999 2210 14033 2239
rect 13999 2142 14033 2166
rect 13999 2074 14033 2092
rect 13999 2006 14033 2018
rect 13999 1938 14033 1944
rect 13999 1830 14033 1836
rect 13999 1756 14033 1768
rect 13999 1682 14033 1700
rect 13999 1608 14033 1632
rect 13999 1548 14033 1564
rect 14135 3104 14255 4200
rect 14135 3070 14178 3104
rect 14212 3070 14255 3104
rect 14135 3026 14255 3070
rect 14135 2992 14178 3026
rect 14212 2992 14255 3026
rect 14135 2948 14255 2992
rect 14135 2914 14178 2948
rect 14212 2914 14255 2948
rect 14135 2870 14255 2914
rect 14135 2836 14178 2870
rect 14212 2836 14255 2870
rect 14135 2792 14255 2836
rect 14135 2758 14178 2792
rect 14212 2758 14255 2792
rect 14135 2713 14255 2758
rect 14135 2679 14178 2713
rect 14212 2679 14255 2713
rect 14135 2634 14255 2679
rect 14135 2600 14178 2634
rect 14212 2600 14255 2634
rect 13777 1470 13820 1504
rect 13854 1470 13897 1504
rect 13777 1430 13897 1470
rect 13777 1396 13820 1430
rect 13854 1396 13897 1430
rect 13777 1250 13897 1396
rect 13777 1144 13784 1250
rect 13890 1144 13897 1250
rect 14135 1504 14255 2600
rect 14135 1470 14178 1504
rect 14212 1470 14255 1504
rect 14135 1430 14255 1470
rect 14135 1396 14178 1430
rect 14212 1396 14255 1430
rect 14135 1250 14255 1396
rect 14135 1144 14142 1250
rect 14248 1144 14255 1250
rect 14356 4286 14428 4325
rect 14390 4252 14428 4286
rect 14356 4213 14428 4252
rect 14390 4179 14428 4213
rect 14356 4140 14428 4179
rect 14390 4106 14428 4140
rect 14356 4082 14428 4106
rect 14390 4033 14428 4082
rect 14356 4014 14428 4033
rect 14390 3960 14428 4014
rect 14356 3957 14536 3960
rect 14356 3952 14468 3957
rect 14356 3946 14428 3952
rect 14390 3918 14428 3946
rect 14462 3923 14468 3952
rect 14502 3924 14536 3957
rect 14502 3923 14604 3924
rect 14462 3921 14604 3923
rect 14462 3918 14500 3921
rect 14390 3888 14500 3918
rect 14534 3889 14572 3921
rect 14638 3905 14653 4551
rect 14390 3887 14468 3888
rect 14534 3887 14536 3889
rect 14356 3880 14468 3887
rect 14356 3878 14428 3880
rect 14390 3846 14428 3878
rect 14462 3854 14468 3880
rect 14502 3855 14536 3887
rect 14570 3887 14572 3889
rect 14606 3887 14653 3905
rect 14570 3871 14653 3887
rect 14570 3855 14604 3871
rect 14502 3854 14604 3855
rect 14462 3848 14604 3854
rect 14462 3846 14500 3848
rect 14390 3819 14500 3846
rect 14534 3820 14572 3848
rect 14638 3837 14653 3871
rect 14390 3814 14468 3819
rect 14534 3814 14536 3820
rect 14356 3810 14468 3814
rect 14390 3808 14468 3810
rect 14390 3776 14428 3808
rect 14356 3775 14428 3776
rect 14390 3774 14428 3775
rect 14462 3785 14468 3808
rect 14502 3786 14536 3814
rect 14570 3814 14572 3820
rect 14606 3814 14653 3837
rect 14570 3803 14653 3814
rect 14570 3786 14604 3803
rect 14502 3785 14604 3786
rect 14462 3775 14604 3785
rect 14462 3774 14500 3775
rect 14390 3750 14500 3774
rect 14534 3751 14572 3775
rect 14638 3769 14653 3803
rect 14390 3736 14468 3750
rect 14534 3741 14536 3751
rect 14390 3708 14428 3736
rect 14356 3702 14428 3708
rect 14462 3716 14468 3736
rect 14502 3717 14536 3741
rect 14570 3741 14572 3751
rect 14606 3741 14653 3769
rect 14570 3735 14653 3741
rect 14570 3717 14604 3735
rect 14502 3716 14604 3717
rect 14462 3702 14604 3716
rect 14390 3681 14500 3702
rect 14534 3682 14572 3702
rect 14638 3701 14653 3735
rect 14390 3664 14468 3681
rect 14534 3668 14536 3682
rect 14390 3640 14428 3664
rect 14356 3630 14428 3640
rect 14462 3647 14468 3664
rect 14502 3648 14536 3668
rect 14570 3668 14572 3682
rect 14606 3668 14653 3701
rect 14570 3667 14653 3668
rect 14570 3648 14604 3667
rect 14502 3647 14604 3648
rect 14462 3633 14604 3647
rect 14638 3633 14653 3667
rect 14462 3630 14653 3633
rect 14356 3629 14653 3630
rect 14390 3612 14500 3629
rect 14534 3613 14572 3629
rect 14390 3592 14468 3612
rect 14534 3595 14536 3613
rect 14390 3572 14428 3592
rect 14356 3558 14428 3572
rect 14462 3578 14468 3592
rect 14502 3579 14536 3595
rect 14570 3595 14572 3613
rect 14606 3599 14653 3629
rect 14570 3579 14604 3595
rect 14502 3578 14604 3579
rect 14462 3565 14604 3578
rect 14638 3565 14653 3599
rect 14462 3558 14653 3565
rect 14356 3556 14653 3558
rect 14390 3543 14500 3556
rect 14534 3544 14572 3556
rect 14390 3520 14468 3543
rect 14534 3522 14536 3544
rect 14390 3504 14428 3520
rect 14356 3486 14428 3504
rect 14462 3509 14468 3520
rect 14502 3510 14536 3522
rect 14570 3522 14572 3544
rect 14606 3531 14653 3556
rect 14570 3510 14604 3522
rect 14502 3509 14604 3510
rect 14462 3497 14604 3509
rect 14638 3497 14653 3531
rect 14462 3486 14653 3497
rect 14356 3483 14653 3486
rect 14390 3474 14500 3483
rect 14534 3475 14572 3483
rect 14390 3448 14468 3474
rect 14534 3449 14536 3475
rect 14390 3436 14428 3448
rect 14356 3414 14428 3436
rect 14462 3440 14468 3448
rect 14502 3441 14536 3449
rect 14570 3449 14572 3475
rect 14606 3463 14653 3483
rect 14570 3441 14604 3449
rect 14502 3440 14604 3441
rect 14462 3429 14604 3440
rect 14638 3429 14653 3463
rect 14462 3414 14653 3429
rect 14356 3410 14653 3414
rect 14390 3405 14500 3410
rect 14534 3406 14572 3410
rect 14390 3376 14468 3405
rect 14534 3376 14536 3406
rect 14390 3368 14428 3376
rect 14356 3342 14428 3368
rect 14462 3371 14468 3376
rect 14502 3372 14536 3376
rect 14570 3376 14572 3406
rect 14606 3395 14653 3410
rect 14570 3372 14604 3376
rect 14502 3371 14604 3372
rect 14462 3361 14604 3371
rect 14638 3361 14653 3395
rect 14462 3342 14653 3361
rect 14356 3337 14653 3342
rect 14390 3336 14500 3337
rect 14390 3304 14468 3336
rect 14390 3300 14428 3304
rect 14356 3270 14428 3300
rect 14462 3302 14468 3304
rect 14534 3303 14536 3337
rect 14570 3303 14572 3337
rect 14606 3327 14653 3337
rect 14502 3302 14604 3303
rect 14462 3293 14604 3302
rect 14638 3293 14653 3327
rect 14462 3270 14653 3293
rect 14356 3268 14653 3270
rect 14356 3267 14536 3268
rect 14356 3266 14468 3267
rect 14390 3233 14468 3266
rect 14502 3264 14536 3267
rect 14534 3234 14536 3264
rect 14570 3264 14653 3268
rect 14570 3234 14572 3264
rect 14606 3259 14653 3264
rect 14390 3232 14500 3233
rect 14390 3230 14428 3232
rect 14356 3198 14428 3230
rect 14462 3230 14500 3232
rect 14534 3230 14572 3234
rect 14462 3225 14604 3230
rect 14638 3225 14653 3259
rect 14462 3199 14653 3225
rect 14462 3198 14536 3199
rect 14390 3164 14468 3198
rect 14502 3191 14536 3198
rect 14534 3165 14536 3191
rect 14570 3191 14653 3199
rect 14570 3165 14572 3191
rect 14390 3160 14500 3164
rect 14390 3157 14428 3160
rect 14356 3126 14428 3157
rect 14462 3157 14500 3160
rect 14534 3157 14572 3165
rect 14638 3157 14653 3191
rect 14462 3130 14653 3157
rect 14462 3129 14536 3130
rect 14462 3126 14468 3129
rect 14356 3118 14468 3126
rect 14502 3118 14536 3129
rect 14390 3095 14468 3118
rect 14534 3096 14536 3118
rect 14570 3123 14653 3130
rect 14570 3118 14604 3123
rect 14570 3096 14572 3118
rect 14390 3088 14500 3095
rect 14390 3084 14428 3088
rect 14356 3054 14428 3084
rect 14462 3084 14500 3088
rect 14534 3084 14572 3096
rect 14638 3089 14653 3123
rect 14606 3084 14653 3089
rect 14462 3061 14653 3084
rect 14462 3060 14536 3061
rect 14462 3054 14468 3060
rect 14356 3045 14468 3054
rect 14502 3045 14536 3060
rect 14390 3026 14468 3045
rect 14534 3027 14536 3045
rect 14570 3055 14653 3061
rect 14570 3045 14604 3055
rect 14570 3027 14572 3045
rect 14390 3016 14500 3026
rect 14390 3011 14428 3016
rect 14356 2982 14428 3011
rect 14462 3011 14500 3016
rect 14534 3011 14572 3027
rect 14638 3021 14653 3055
rect 14606 3011 14653 3021
rect 14462 2992 14653 3011
rect 14462 2991 14536 2992
rect 14462 2982 14468 2991
rect 14356 2972 14468 2982
rect 14502 2972 14536 2991
rect 14390 2957 14468 2972
rect 14534 2958 14536 2972
rect 14570 2987 14653 2992
rect 14570 2972 14604 2987
rect 14570 2958 14572 2972
rect 14390 2944 14500 2957
rect 14390 2938 14428 2944
rect 14356 2910 14428 2938
rect 14462 2938 14500 2944
rect 14534 2938 14572 2958
rect 14638 2953 14653 2987
rect 14606 2938 14653 2953
rect 14462 2923 14653 2938
rect 14462 2922 14536 2923
rect 14462 2910 14468 2922
rect 14356 2899 14468 2910
rect 14502 2899 14536 2922
rect 14390 2888 14468 2899
rect 14534 2889 14536 2899
rect 14570 2919 14653 2923
rect 14570 2899 14604 2919
rect 14570 2889 14572 2899
rect 14390 2872 14500 2888
rect 14390 2865 14428 2872
rect 14356 2838 14428 2865
rect 14462 2865 14500 2872
rect 14534 2865 14572 2889
rect 14638 2885 14653 2919
rect 14606 2865 14653 2885
rect 14462 2854 14653 2865
rect 14462 2853 14536 2854
rect 14462 2838 14468 2853
rect 14356 2826 14468 2838
rect 14502 2826 14536 2853
rect 14390 2819 14468 2826
rect 14534 2820 14536 2826
rect 14570 2851 14653 2854
rect 14570 2826 14604 2851
rect 14570 2820 14572 2826
rect 14390 2800 14500 2819
rect 14390 2792 14428 2800
rect 14356 2766 14428 2792
rect 14462 2792 14500 2800
rect 14534 2792 14572 2820
rect 14638 2817 14653 2851
rect 14606 2792 14653 2817
rect 14462 2785 14653 2792
rect 14462 2784 14536 2785
rect 14462 2766 14468 2784
rect 14356 2753 14468 2766
rect 14502 2753 14536 2784
rect 14390 2750 14468 2753
rect 14534 2751 14536 2753
rect 14570 2783 14653 2785
rect 14570 2753 14604 2783
rect 14570 2751 14572 2753
rect 14390 2728 14500 2750
rect 14390 2719 14428 2728
rect 14356 2694 14428 2719
rect 14462 2719 14500 2728
rect 14534 2719 14572 2751
rect 14638 2749 14653 2783
rect 14606 2719 14653 2749
rect 14462 2716 14653 2719
rect 14462 2715 14536 2716
rect 14462 2694 14468 2715
rect 14356 2681 14468 2694
rect 14502 2682 14536 2715
rect 14570 2715 14653 2716
rect 14570 2682 14604 2715
rect 14502 2681 14604 2682
rect 14638 2681 14653 2715
rect 14356 2680 14653 2681
rect 14390 2656 14500 2680
rect 14390 2646 14428 2656
rect 14356 2622 14428 2646
rect 14462 2646 14500 2656
rect 14534 2647 14572 2680
rect 14606 2647 14653 2680
rect 14534 2646 14536 2647
rect 14462 2622 14468 2646
rect 14356 2612 14468 2622
rect 14502 2613 14536 2646
rect 14570 2646 14572 2647
rect 14570 2613 14604 2646
rect 14638 2613 14653 2647
rect 14502 2612 14653 2613
rect 14356 2607 14653 2612
rect 14390 2584 14500 2607
rect 14390 2573 14428 2584
rect 14356 2550 14428 2573
rect 14462 2577 14500 2584
rect 14534 2578 14572 2607
rect 14606 2579 14653 2607
rect 14462 2550 14468 2577
rect 14534 2573 14536 2578
rect 14356 2543 14468 2550
rect 14502 2544 14536 2573
rect 14570 2573 14572 2578
rect 14570 2545 14604 2573
rect 14638 2545 14653 2579
rect 14570 2544 14653 2545
rect 14502 2543 14653 2544
rect 14356 2534 14653 2543
rect 14390 2512 14500 2534
rect 14390 2500 14428 2512
rect 14356 2482 14428 2500
rect 14390 2478 14428 2482
rect 14462 2508 14500 2512
rect 14534 2509 14572 2534
rect 14606 2511 14653 2534
rect 14462 2478 14468 2508
rect 14534 2500 14536 2509
rect 14390 2474 14468 2478
rect 14502 2475 14536 2500
rect 14570 2500 14572 2509
rect 14570 2477 14604 2500
rect 14638 2477 14653 2511
rect 14570 2475 14653 2477
rect 14502 2474 14653 2475
rect 14390 2461 14653 2474
rect 14390 2440 14500 2461
rect 14390 2427 14428 2440
rect 14356 2414 14428 2427
rect 14390 2406 14428 2414
rect 14462 2439 14500 2440
rect 14534 2440 14572 2461
rect 14606 2443 14653 2461
rect 14462 2406 14468 2439
rect 14534 2427 14536 2440
rect 14390 2405 14468 2406
rect 14502 2406 14536 2427
rect 14570 2427 14572 2440
rect 14570 2409 14604 2427
rect 14638 2409 14653 2443
rect 14570 2406 14653 2409
rect 14502 2405 14653 2406
rect 14390 2388 14653 2405
rect 14390 2370 14500 2388
rect 14534 2371 14572 2388
rect 14606 2375 14653 2388
rect 14390 2368 14468 2370
rect 14390 2354 14428 2368
rect 14356 2346 14428 2354
rect 14390 2334 14428 2346
rect 14462 2336 14468 2368
rect 14534 2354 14536 2371
rect 14502 2337 14536 2354
rect 14570 2354 14572 2371
rect 14570 2341 14604 2354
rect 14638 2341 14653 2375
rect 14570 2337 14653 2341
rect 14502 2336 14653 2337
rect 14462 2334 14653 2336
rect 14390 2315 14653 2334
rect 14390 2301 14500 2315
rect 14534 2302 14572 2315
rect 14606 2307 14653 2315
rect 14390 2296 14468 2301
rect 14390 2281 14428 2296
rect 14356 2278 14428 2281
rect 14390 2262 14428 2278
rect 14462 2267 14468 2296
rect 14534 2281 14536 2302
rect 14502 2268 14536 2281
rect 14570 2281 14572 2302
rect 14570 2273 14604 2281
rect 14638 2273 14653 2307
rect 14570 2268 14653 2273
rect 14502 2267 14653 2268
rect 14462 2262 14653 2267
rect 14390 2244 14653 2262
rect 14356 2242 14653 2244
rect 14390 2232 14500 2242
rect 14534 2233 14572 2242
rect 14606 2239 14653 2242
rect 14390 2224 14468 2232
rect 14390 2190 14428 2224
rect 14462 2198 14468 2224
rect 14534 2208 14536 2233
rect 14502 2199 14536 2208
rect 14570 2208 14572 2233
rect 14570 2205 14604 2208
rect 14638 2205 14653 2239
rect 14570 2199 14653 2205
rect 14502 2198 14653 2199
rect 14462 2190 14653 2198
rect 14390 2176 14653 2190
rect 14356 2171 14653 2176
rect 14356 2169 14604 2171
rect 14390 2163 14500 2169
rect 14534 2164 14572 2169
rect 14390 2152 14468 2163
rect 14390 2118 14428 2152
rect 14462 2129 14468 2152
rect 14534 2135 14536 2164
rect 14502 2130 14536 2135
rect 14570 2135 14572 2164
rect 14638 2137 14653 2171
rect 14606 2135 14653 2137
rect 14570 2130 14653 2135
rect 14502 2129 14653 2130
rect 14462 2118 14653 2129
rect 14390 2108 14653 2118
rect 14356 2103 14653 2108
rect 14356 2096 14604 2103
rect 14390 2094 14500 2096
rect 14534 2095 14572 2096
rect 14390 2080 14468 2094
rect 14390 2046 14428 2080
rect 14462 2060 14468 2080
rect 14534 2062 14536 2095
rect 14502 2061 14536 2062
rect 14570 2062 14572 2095
rect 14638 2069 14653 2103
rect 14606 2062 14653 2069
rect 14570 2061 14653 2062
rect 14502 2060 14653 2061
rect 14462 2046 14653 2060
rect 14390 2040 14653 2046
rect 14356 2035 14653 2040
rect 14356 2026 14604 2035
rect 14356 2025 14536 2026
rect 14356 2023 14468 2025
rect 14502 2023 14536 2025
rect 14390 2008 14468 2023
rect 14390 1974 14428 2008
rect 14462 1991 14468 2008
rect 14534 1992 14536 2023
rect 14570 2023 14604 2026
rect 14570 1992 14572 2023
rect 14638 2001 14653 2035
rect 14462 1989 14500 1991
rect 14534 1989 14572 1992
rect 14606 1989 14653 2001
rect 14462 1974 14653 1989
rect 14390 1972 14653 1974
rect 14356 1967 14653 1972
rect 14356 1957 14604 1967
rect 14356 1956 14536 1957
rect 14356 1950 14468 1956
rect 14502 1950 14536 1956
rect 14390 1936 14468 1950
rect 14390 1904 14428 1936
rect 14356 1902 14428 1904
rect 14462 1922 14468 1936
rect 14534 1923 14536 1950
rect 14570 1950 14604 1957
rect 14570 1923 14572 1950
rect 14638 1933 14653 1967
rect 14462 1916 14500 1922
rect 14534 1916 14572 1923
rect 14606 1916 14653 1933
rect 14462 1902 14653 1916
rect 14356 1899 14653 1902
rect 14356 1888 14604 1899
rect 14356 1887 14536 1888
rect 14356 1877 14468 1887
rect 14502 1877 14536 1887
rect 14390 1864 14468 1877
rect 14390 1836 14428 1864
rect 14356 1830 14428 1836
rect 14462 1853 14468 1864
rect 14534 1854 14536 1877
rect 14570 1877 14604 1888
rect 14570 1854 14572 1877
rect 14638 1865 14653 1899
rect 14462 1843 14500 1853
rect 14534 1843 14572 1854
rect 14606 1843 14653 1865
rect 14462 1831 14653 1843
rect 14462 1830 14604 1831
rect 14356 1819 14604 1830
rect 14356 1818 14536 1819
rect 14356 1804 14468 1818
rect 14502 1804 14536 1818
rect 14390 1792 14468 1804
rect 14390 1768 14428 1792
rect 14356 1758 14428 1768
rect 14462 1784 14468 1792
rect 14534 1785 14536 1804
rect 14570 1804 14604 1819
rect 14570 1785 14572 1804
rect 14638 1797 14653 1831
rect 14462 1770 14500 1784
rect 14534 1770 14572 1785
rect 14606 1770 14653 1797
rect 14462 1763 14653 1770
rect 14462 1758 14604 1763
rect 14356 1750 14604 1758
rect 14356 1749 14536 1750
rect 14356 1734 14468 1749
rect 14390 1720 14468 1734
rect 14502 1731 14536 1749
rect 14390 1697 14428 1720
rect 14356 1686 14428 1697
rect 14462 1715 14468 1720
rect 14534 1716 14536 1731
rect 14570 1731 14604 1750
rect 14570 1716 14572 1731
rect 14638 1729 14653 1763
rect 14462 1697 14500 1715
rect 14534 1697 14572 1716
rect 14606 1697 14653 1729
rect 14462 1695 14653 1697
rect 14462 1686 14604 1695
rect 14356 1681 14604 1686
rect 14356 1680 14536 1681
rect 14356 1666 14468 1680
rect 14390 1648 14468 1666
rect 14502 1658 14536 1680
rect 14390 1623 14428 1648
rect 14356 1614 14428 1623
rect 14462 1646 14468 1648
rect 14534 1647 14536 1658
rect 14570 1661 14604 1681
rect 14638 1661 14653 1695
rect 14570 1658 14653 1661
rect 14570 1647 14572 1658
rect 14462 1624 14500 1646
rect 14534 1624 14572 1647
rect 14606 1627 14653 1658
rect 14462 1614 14604 1624
rect 14356 1612 14604 1614
rect 14356 1611 14536 1612
rect 14356 1598 14468 1611
rect 14390 1577 14468 1598
rect 14502 1585 14536 1611
rect 14534 1578 14536 1585
rect 14570 1593 14604 1612
rect 14638 1593 14653 1627
rect 14570 1585 14653 1593
rect 14570 1578 14572 1585
rect 14390 1576 14500 1577
rect 14390 1549 14428 1576
rect 14356 1542 14428 1549
rect 14462 1551 14500 1576
rect 14534 1551 14572 1578
rect 14606 1559 14653 1585
rect 14462 1543 14604 1551
rect 14462 1542 14536 1543
rect 14356 1509 14468 1542
rect 14502 1512 14536 1542
rect 14390 1508 14468 1509
rect 14534 1509 14536 1512
rect 14570 1525 14604 1543
rect 14638 1525 14653 1559
rect 14570 1512 14653 1525
rect 14570 1509 14572 1512
rect 14390 1504 14500 1508
rect 14390 1475 14428 1504
rect 14356 1470 14428 1475
rect 14462 1478 14500 1504
rect 14534 1478 14572 1509
rect 14606 1491 14653 1512
rect 14462 1474 14604 1478
rect 14462 1473 14536 1474
rect 14462 1470 14468 1473
rect 14356 1439 14468 1470
rect 14502 1440 14536 1473
rect 14570 1457 14604 1474
rect 14638 1457 14653 1491
rect 14570 1440 14653 1457
rect 14502 1439 14653 1440
rect 14356 1435 14500 1439
rect 14390 1432 14500 1435
rect 14390 1401 14428 1432
rect 14356 1398 14428 1401
rect 14462 1405 14500 1432
rect 14534 1405 14572 1439
rect 14606 1423 14653 1439
rect 14462 1404 14536 1405
rect 14462 1398 14468 1404
rect 14356 1370 14468 1398
rect 14502 1371 14536 1404
rect 14570 1389 14604 1405
rect 14638 1389 14653 1423
rect 14570 1371 14653 1389
rect 14502 1370 14653 1371
rect 14356 1366 14653 1370
rect 14356 1361 14500 1366
rect 14390 1360 14500 1361
rect 14390 1327 14428 1360
rect 14356 1326 14428 1327
rect 14462 1335 14500 1360
rect 14534 1336 14572 1366
rect 14606 1355 14653 1366
rect 14462 1326 14468 1335
rect 14534 1332 14536 1336
rect 14356 1301 14468 1326
rect 14502 1302 14536 1332
rect 14570 1332 14572 1336
rect 14570 1321 14604 1332
rect 14638 1321 14653 1355
rect 14570 1302 14653 1321
rect 14502 1301 14653 1302
rect 14356 1293 14653 1301
rect 14356 1288 14500 1293
rect 14356 1287 14428 1288
rect 14390 1254 14428 1287
rect 14462 1266 14500 1288
rect 14534 1267 14572 1293
rect 14606 1287 14653 1293
rect 14462 1254 14468 1266
rect 14534 1259 14536 1267
rect 14390 1253 14468 1254
rect 14356 1232 14468 1253
rect 14502 1233 14536 1259
rect 14570 1259 14572 1267
rect 14570 1253 14604 1259
rect 14638 1253 14653 1287
rect 14570 1233 14653 1253
rect 14502 1232 14653 1233
rect 14356 1220 14653 1232
rect 14356 1216 14500 1220
rect 14356 1213 14428 1216
rect 14390 1182 14428 1213
rect 14462 1197 14500 1216
rect 14534 1198 14572 1220
rect 14606 1218 14653 1220
rect 14462 1182 14468 1197
rect 14534 1186 14536 1198
rect 14390 1179 14468 1182
rect 14356 1163 14468 1179
rect 14502 1164 14536 1186
rect 14570 1186 14572 1198
rect 14570 1184 14604 1186
rect 14638 1184 14653 1218
rect 14570 1164 14653 1184
rect 14502 1163 14653 1164
rect 14356 1149 14653 1163
rect 14356 1147 14604 1149
rect 14356 1144 14500 1147
rect 667 883 746 894
rect 667 867 780 883
rect 14356 1139 14428 1144
rect 14390 1110 14428 1139
rect 14462 1128 14500 1144
rect 14534 1129 14572 1147
rect 14462 1110 14468 1128
rect 14534 1113 14536 1129
rect 14390 1105 14468 1110
rect 14356 1094 14468 1105
rect 14502 1095 14536 1113
rect 14570 1113 14572 1129
rect 14638 1115 14653 1149
rect 14606 1113 14653 1115
rect 14570 1095 14653 1113
rect 14502 1094 14653 1095
rect 14356 1080 14653 1094
rect 14356 1074 14604 1080
rect 14356 1072 14500 1074
rect 14356 1065 14428 1072
rect 14390 1038 14428 1065
rect 14462 1059 14500 1072
rect 14534 1060 14572 1074
rect 14462 1038 14468 1059
rect 14534 1040 14536 1060
rect 14390 1031 14468 1038
rect 14356 1025 14468 1031
rect 14502 1026 14536 1040
rect 14570 1040 14572 1060
rect 14638 1046 14653 1080
rect 14606 1040 14653 1046
rect 14570 1026 14653 1040
rect 14502 1025 14653 1026
rect 14356 1011 14653 1025
rect 14356 1001 14604 1011
rect 14356 1000 14500 1001
rect 14356 991 14428 1000
rect 14390 966 14428 991
rect 14462 990 14500 1000
rect 14534 991 14572 1001
rect 14462 966 14468 990
rect 14534 967 14536 991
rect 14390 957 14468 966
rect 14356 956 14468 957
rect 14502 957 14536 967
rect 14570 967 14572 991
rect 14638 977 14653 1011
rect 14606 967 14653 977
rect 14570 957 14653 967
rect 14502 956 14653 957
rect 14356 942 14653 956
rect 14356 928 14604 942
rect 14356 917 14428 928
rect 14390 894 14428 917
rect 14462 921 14500 928
rect 14534 922 14572 928
rect 14462 894 14468 921
rect 14534 894 14536 922
rect 14390 887 14468 894
rect 14502 888 14536 894
rect 14570 894 14572 922
rect 14638 908 14653 942
rect 14606 894 14653 908
rect 14570 888 14653 894
rect 14502 887 14653 888
rect 14390 883 14653 887
rect 14356 873 14653 883
rect 14356 867 14604 873
rect 667 853 14604 867
rect 667 852 14536 853
rect 667 818 702 852
rect 736 820 771 852
rect 805 820 840 852
rect 874 820 909 852
rect 943 820 978 852
rect 1012 820 1047 852
rect 1081 820 1116 852
rect 1150 820 1185 852
rect 1219 820 1254 852
rect 1288 820 1323 852
rect 1357 820 1392 852
rect 1426 820 1461 852
rect 1495 820 1530 852
rect 1564 820 1599 852
rect 1633 820 1668 852
rect 1702 820 1737 852
rect 1771 820 1806 852
rect 1840 820 1875 852
rect 1909 820 1944 852
rect 1978 820 2013 852
rect 2047 820 2082 852
rect 2116 820 2151 852
rect 2185 820 2220 852
rect 2254 820 2289 852
rect 2323 820 2358 852
rect 2392 820 2427 852
rect 2461 820 2496 852
rect 2530 820 2565 852
rect 2599 820 2634 852
rect 2668 820 2703 852
rect 2737 820 2772 852
rect 743 818 771 820
rect 816 818 840 820
rect 889 818 909 820
rect 599 786 709 818
rect 743 786 782 818
rect 816 786 855 818
rect 889 786 928 818
rect 599 784 928 786
rect 482 750 565 769
rect 599 750 634 784
rect 668 750 703 784
rect 737 750 772 784
rect 806 750 841 784
rect 875 750 910 784
rect 14502 819 14536 852
rect 14570 839 14604 853
rect 14638 839 14653 873
rect 14570 819 14653 839
rect 14502 804 14653 819
rect 14502 784 14604 804
rect 14570 770 14604 784
rect 14638 770 14653 804
rect 14570 750 14653 770
rect 482 748 928 750
rect 482 716 709 748
rect 743 716 782 748
rect 816 716 855 748
rect 889 716 928 748
rect 482 682 516 716
rect 550 682 585 716
rect 619 682 654 716
rect 688 714 709 716
rect 757 714 782 716
rect 826 714 855 716
rect 895 714 928 716
rect 14551 735 14653 750
rect 688 682 723 714
rect 757 682 792 714
rect 826 682 861 714
rect 895 682 930 714
rect 964 682 999 714
rect 1033 682 1068 714
rect 1102 682 1137 714
rect 1171 682 1206 714
rect 1240 682 1275 714
rect 1309 682 1344 714
rect 1378 682 1413 714
rect 1447 682 1482 714
rect 1516 682 1551 714
rect 1585 682 1620 714
rect 1654 682 1689 714
rect 1723 682 1758 714
rect 1792 682 1827 714
rect 1861 682 1896 714
rect 1930 682 1965 714
rect 1999 682 2034 714
rect 2068 682 2103 714
rect 2137 682 2172 714
rect 2206 682 2241 714
rect 2275 682 2310 714
rect 2344 682 2379 714
rect 2413 682 2448 714
rect 2482 682 2517 714
rect 2551 682 2586 714
rect 2620 682 2655 714
rect 2689 682 2724 714
rect 2758 682 2793 714
rect 2827 682 2862 714
rect 2896 682 2931 714
rect 2965 682 3000 714
rect 3034 682 3069 714
rect 3103 682 3138 714
rect 3172 682 3207 714
rect 3241 682 3276 714
rect 3310 682 3345 714
rect 3379 682 3414 714
rect 3448 682 3483 714
rect 3517 682 3552 714
rect 3586 682 3621 714
rect 3655 682 3690 714
rect 3724 682 3759 714
rect 3793 682 3828 714
rect 3862 682 3897 714
rect 3931 682 3966 714
rect 4000 682 4035 714
rect 4069 682 4104 714
rect 4138 682 4173 714
rect 4207 682 4242 714
rect 4276 682 4311 714
rect 4345 682 4380 714
rect 4414 682 4449 714
rect 4483 682 4518 714
rect 4552 682 4587 714
rect 4621 682 4656 714
rect 4690 682 4725 714
rect 14551 701 14604 735
rect 14638 701 14653 735
rect 14551 682 14653 701
rect 482 667 14653 682
rect 14807 4636 14832 4670
rect 14866 4655 14907 4670
rect 14807 4621 14840 4636
rect 14874 4621 14907 4655
rect 14807 4598 14907 4621
rect 14807 4564 14832 4598
rect 14866 4587 14907 4598
rect 14807 4553 14840 4564
rect 14874 4553 14907 4587
rect 14807 4526 14907 4553
rect 14807 4492 14832 4526
rect 14866 4519 14907 4526
rect 14807 4485 14840 4492
rect 14874 4485 14907 4519
rect 14807 4454 14907 4485
rect 14807 4420 14832 4454
rect 14866 4451 14907 4454
rect 14807 4417 14840 4420
rect 14874 4417 14907 4451
rect 14807 4383 14907 4417
rect 14807 4382 14840 4383
rect 14807 4348 14832 4382
rect 14874 4349 14907 4383
rect 14866 4348 14907 4349
rect 14807 4315 14907 4348
rect 14807 4310 14840 4315
rect 14807 4276 14832 4310
rect 14874 4281 14907 4315
rect 14866 4276 14907 4281
rect 14807 4247 14907 4276
rect 14807 4238 14840 4247
rect 14807 4204 14832 4238
rect 14874 4213 14907 4247
rect 14866 4204 14907 4213
rect 14807 4179 14907 4204
rect 14807 4166 14840 4179
rect 14807 4132 14832 4166
rect 14874 4145 14907 4179
rect 14866 4132 14907 4145
rect 14807 4111 14907 4132
rect 14807 4094 14840 4111
rect 14807 4060 14832 4094
rect 14874 4077 14907 4111
rect 14866 4060 14907 4077
rect 14807 4043 14907 4060
rect 14807 4022 14840 4043
rect 14807 3988 14832 4022
rect 14874 4009 14907 4043
rect 14866 3988 14907 4009
rect 14807 3975 14907 3988
rect 14807 3950 14840 3975
rect 14807 3916 14832 3950
rect 14874 3941 14907 3975
rect 14866 3916 14907 3941
rect 14807 3907 14907 3916
rect 14807 3878 14840 3907
rect 14807 3844 14832 3878
rect 14874 3873 14907 3907
rect 14866 3844 14907 3873
rect 14807 3839 14907 3844
rect 14807 3806 14840 3839
rect 14807 3772 14832 3806
rect 14874 3805 14907 3839
rect 14866 3772 14907 3805
rect 14807 3771 14907 3772
rect 14807 3737 14840 3771
rect 14874 3737 14907 3771
rect 14807 3734 14907 3737
rect 14807 3700 14832 3734
rect 14866 3703 14907 3734
rect 14807 3669 14840 3700
rect 14874 3669 14907 3703
rect 14807 3662 14907 3669
rect 14807 3628 14832 3662
rect 14866 3635 14907 3662
rect 14807 3601 14840 3628
rect 14874 3601 14907 3635
rect 14807 3590 14907 3601
rect 14807 3556 14832 3590
rect 14866 3567 14907 3590
rect 14807 3533 14840 3556
rect 14874 3533 14907 3567
rect 14807 3518 14907 3533
rect 14807 3484 14832 3518
rect 14866 3499 14907 3518
rect 14807 3465 14840 3484
rect 14874 3465 14907 3499
rect 14807 3446 14907 3465
rect 14807 3412 14832 3446
rect 14866 3431 14907 3446
rect 14807 3397 14840 3412
rect 14874 3397 14907 3431
rect 14807 3374 14907 3397
rect 14807 3340 14832 3374
rect 14866 3363 14907 3374
rect 14807 3329 14840 3340
rect 14874 3329 14907 3363
rect 14807 3302 14907 3329
rect 14807 3268 14832 3302
rect 14866 3295 14907 3302
rect 14807 3261 14840 3268
rect 14874 3261 14907 3295
rect 14807 3230 14907 3261
rect 14807 3196 14832 3230
rect 14866 3227 14907 3230
rect 14807 3193 14840 3196
rect 14874 3193 14907 3227
rect 14807 3159 14907 3193
rect 14807 3158 14840 3159
rect 14807 3124 14832 3158
rect 14874 3125 14907 3159
rect 14866 3124 14907 3125
rect 14807 3091 14907 3124
rect 14807 3086 14840 3091
rect 14807 3052 14832 3086
rect 14874 3057 14907 3091
rect 14866 3052 14907 3057
rect 14807 3023 14907 3052
rect 14807 3014 14840 3023
rect 14807 2980 14832 3014
rect 14874 2989 14907 3023
rect 14866 2980 14907 2989
rect 14807 2955 14907 2980
rect 14807 2942 14840 2955
rect 14807 2908 14832 2942
rect 14874 2921 14907 2955
rect 14866 2908 14907 2921
rect 14807 2887 14907 2908
rect 14807 2870 14840 2887
rect 14807 2836 14832 2870
rect 14874 2853 14907 2887
rect 14866 2836 14907 2853
rect 14807 2819 14907 2836
rect 14807 2798 14840 2819
rect 14807 2764 14832 2798
rect 14874 2785 14907 2819
rect 14866 2764 14907 2785
rect 14807 2751 14907 2764
rect 14807 2726 14840 2751
rect 14807 2692 14832 2726
rect 14874 2717 14907 2751
rect 14866 2692 14907 2717
rect 14807 2683 14907 2692
rect 14807 2654 14840 2683
rect 14807 2620 14832 2654
rect 14874 2649 14907 2683
rect 14866 2620 14907 2649
rect 14807 2615 14907 2620
rect 14807 2582 14840 2615
rect 14807 2548 14832 2582
rect 14874 2581 14907 2615
rect 14866 2548 14907 2581
rect 14807 2547 14907 2548
rect 14807 2513 14840 2547
rect 14874 2513 14907 2547
rect 14807 2510 14907 2513
rect 14807 2476 14832 2510
rect 14866 2479 14907 2510
rect 14807 2445 14840 2476
rect 14874 2445 14907 2479
rect 14807 2438 14907 2445
rect 14807 2404 14832 2438
rect 14866 2411 14907 2438
rect 14807 2377 14840 2404
rect 14874 2377 14907 2411
rect 14807 2366 14907 2377
rect 14807 2332 14832 2366
rect 14866 2343 14907 2366
rect 14807 2309 14840 2332
rect 14874 2309 14907 2343
rect 14807 2294 14907 2309
rect 14807 2260 14832 2294
rect 14866 2275 14907 2294
rect 14807 2241 14840 2260
rect 14874 2241 14907 2275
rect 14807 2222 14907 2241
rect 14807 2188 14832 2222
rect 14866 2207 14907 2222
rect 14807 2173 14840 2188
rect 14874 2173 14907 2207
rect 14807 2150 14907 2173
rect 14807 2116 14832 2150
rect 14866 2139 14907 2150
rect 14807 2105 14840 2116
rect 14874 2105 14907 2139
rect 14807 2078 14907 2105
rect 14807 2044 14832 2078
rect 14866 2071 14907 2078
rect 14807 2037 14840 2044
rect 14874 2037 14907 2071
rect 14807 2006 14907 2037
rect 14807 1972 14832 2006
rect 14866 2003 14907 2006
rect 14807 1969 14840 1972
rect 14874 1969 14907 2003
rect 14807 1935 14907 1969
rect 14807 1934 14840 1935
rect 14807 1900 14832 1934
rect 14874 1901 14907 1935
rect 14866 1900 14907 1901
rect 14807 1867 14907 1900
rect 14807 1862 14840 1867
rect 14807 1828 14832 1862
rect 14874 1833 14907 1867
rect 14866 1828 14907 1833
rect 14807 1799 14907 1828
rect 14807 1790 14840 1799
rect 14807 1756 14832 1790
rect 14874 1765 14907 1799
rect 14866 1756 14907 1765
rect 14807 1731 14907 1756
rect 14807 1718 14840 1731
rect 14807 1684 14832 1718
rect 14874 1697 14907 1731
rect 14866 1684 14907 1697
rect 14807 1663 14907 1684
rect 14807 1646 14840 1663
rect 14807 1612 14832 1646
rect 14874 1629 14907 1663
rect 14866 1612 14907 1629
rect 14807 1595 14907 1612
rect 14807 1574 14840 1595
rect 14807 1540 14832 1574
rect 14874 1561 14907 1595
rect 14866 1540 14907 1561
rect 14807 1527 14907 1540
rect 14807 1502 14840 1527
rect 14807 1468 14832 1502
rect 14874 1493 14907 1527
rect 14866 1468 14907 1493
rect 14807 1459 14907 1468
rect 14807 1429 14840 1459
rect 14807 1395 14832 1429
rect 14874 1425 14907 1459
rect 14866 1395 14907 1425
rect 14807 1391 14907 1395
rect 14807 1357 14840 1391
rect 14874 1357 14907 1391
rect 14807 1356 14907 1357
rect 14807 1322 14832 1356
rect 14866 1323 14907 1356
rect 14807 1289 14840 1322
rect 14874 1289 14907 1323
rect 14807 1283 14907 1289
rect 14807 1249 14832 1283
rect 14866 1255 14907 1283
rect 14807 1221 14840 1249
rect 14874 1221 14907 1255
rect 14807 1210 14907 1221
rect 14807 1176 14832 1210
rect 14866 1187 14907 1210
rect 14807 1153 14840 1176
rect 14874 1153 14907 1187
rect 14807 1137 14907 1153
rect 14807 1103 14832 1137
rect 14866 1119 14907 1137
rect 14807 1085 14840 1103
rect 14874 1085 14907 1119
rect 14807 1064 14907 1085
rect 14807 1030 14832 1064
rect 14866 1051 14907 1064
rect 14807 1017 14840 1030
rect 14874 1017 14907 1051
rect 14807 991 14907 1017
rect 14807 957 14832 991
rect 14866 983 14907 991
rect 14807 949 14840 957
rect 14874 949 14907 983
rect 14807 918 14907 949
rect 14807 884 14832 918
rect 14866 915 14907 918
rect 14807 881 14840 884
rect 14874 881 14907 915
rect 14807 847 14907 881
rect 14807 845 14840 847
rect 14807 811 14832 845
rect 14874 813 14907 847
rect 14866 811 14907 813
rect 14807 779 14907 811
rect 14807 772 14840 779
rect 14807 738 14832 772
rect 14874 745 14907 779
rect 14866 738 14907 745
rect 14807 711 14907 738
rect 14807 699 14840 711
rect 229 609 262 643
rect 296 641 329 643
rect 229 607 269 609
rect 303 607 329 641
rect 229 575 329 607
rect 229 541 262 575
rect 296 567 329 575
rect 229 533 269 541
rect 303 533 329 567
rect 229 514 329 533
rect 14807 665 14832 699
rect 14874 677 14907 711
rect 14866 665 14907 677
rect 14807 643 14907 665
rect 14807 626 14840 643
rect 14807 592 14832 626
rect 14874 609 14907 643
rect 14866 592 14907 609
rect 14807 575 14907 592
rect 14807 553 14840 575
rect 14807 519 14832 553
rect 14874 541 14907 575
rect 14866 519 14907 541
rect 14807 514 14907 519
rect 229 499 14907 514
rect 229 465 302 499
rect 336 497 375 499
rect 409 497 448 499
rect 482 497 521 499
rect 555 497 594 499
rect 628 497 667 499
rect 336 465 343 497
rect 409 465 419 497
rect 482 465 495 497
rect 555 465 571 497
rect 628 465 648 497
rect 701 465 740 499
rect 774 465 813 499
rect 847 465 886 499
rect 920 465 959 499
rect 993 465 1032 499
rect 1066 465 1105 499
rect 1139 465 1178 499
rect 1212 465 1251 499
rect 1285 465 1324 499
rect 1358 465 1397 499
rect 1431 465 1470 499
rect 1504 465 1543 499
rect 1577 465 1616 499
rect 1650 465 1689 499
rect 1723 465 1762 499
rect 1796 465 1835 499
rect 1869 465 1908 499
rect 1942 465 1981 499
rect 2015 465 2054 499
rect 2088 465 2127 499
rect 2161 465 2200 499
rect 2234 465 2273 499
rect 2307 465 2346 499
rect 2380 465 2419 499
rect 2453 465 2492 499
rect 2526 465 2565 499
rect 2599 465 2638 499
rect 2672 465 2711 499
rect 2745 465 2784 499
rect 2818 465 2857 499
rect 2891 465 2930 499
rect 2964 465 3003 499
rect 3037 465 3076 499
rect 3110 465 3149 499
rect 3183 465 3222 499
rect 3256 465 3295 499
rect 3329 465 3368 499
rect 3402 465 3441 499
rect 3475 465 3514 499
rect 3548 465 3587 499
rect 3621 465 3660 499
rect 3694 465 3733 499
rect 3767 465 3806 499
rect 3840 465 3879 499
rect 3913 465 3952 499
rect 3986 465 4025 499
rect 4059 465 4098 499
rect 4132 465 4171 499
rect 4205 465 4244 499
rect 4278 465 4317 499
rect 4351 465 4390 499
rect 4424 465 4463 499
rect 4497 465 4536 499
rect 4570 465 4609 499
rect 4643 465 4682 499
rect 4716 465 4755 499
rect 4789 465 4828 499
rect 4862 465 4901 499
rect 4935 465 4974 499
rect 5008 465 5047 499
rect 5081 465 5120 499
rect 5154 465 5193 499
rect 5227 465 5266 499
rect 5300 465 5339 499
rect 5373 465 5411 499
rect 5445 465 5483 499
rect 5517 465 5555 499
rect 5589 465 5627 499
rect 5661 465 5699 499
rect 5733 465 5771 499
rect 5805 465 5843 499
rect 5877 465 5915 499
rect 5949 465 5987 499
rect 6021 465 6059 499
rect 6093 465 6131 499
rect 6165 465 6203 499
rect 6237 465 6275 499
rect 6309 465 6347 499
rect 6381 465 6419 499
rect 6453 465 6491 499
rect 6525 465 6563 499
rect 6597 465 6635 499
rect 6669 465 6707 499
rect 6741 465 6779 499
rect 6813 465 6851 499
rect 6885 465 6923 499
rect 6957 465 6995 499
rect 7029 465 7067 499
rect 7101 465 7139 499
rect 7173 465 7211 499
rect 7245 465 7283 499
rect 7317 465 7355 499
rect 7389 465 7427 499
rect 7461 465 7499 499
rect 7533 465 7571 499
rect 7605 465 7643 499
rect 7677 465 7715 499
rect 7749 465 7787 499
rect 7821 465 7859 499
rect 7893 465 7931 499
rect 7965 465 8003 499
rect 8037 465 8075 499
rect 8109 465 8147 499
rect 8181 465 8219 499
rect 8253 465 8291 499
rect 8325 465 8363 499
rect 8397 465 8435 499
rect 8469 465 8507 499
rect 8541 465 8579 499
rect 8613 465 8651 499
rect 8685 465 8723 499
rect 8757 465 8795 499
rect 8829 465 8867 499
rect 8901 465 8939 499
rect 8973 465 9011 499
rect 9045 465 9083 499
rect 9117 465 9155 499
rect 9189 465 9227 499
rect 9261 465 9299 499
rect 9333 465 9371 499
rect 9405 465 9443 499
rect 9477 465 9515 499
rect 9549 465 9587 499
rect 9621 465 9659 499
rect 9693 465 9731 499
rect 9765 465 9803 499
rect 9837 465 9875 499
rect 9909 465 9947 499
rect 9981 465 10019 499
rect 10053 465 10091 499
rect 10125 465 10163 499
rect 10197 465 10235 499
rect 10269 465 10307 499
rect 10341 465 10379 499
rect 10413 465 10451 499
rect 10485 465 10523 499
rect 10557 465 10595 499
rect 10629 465 10667 499
rect 10701 465 10739 499
rect 10773 465 10811 499
rect 10845 465 10883 499
rect 10917 465 10955 499
rect 10989 465 11027 499
rect 11061 465 11099 499
rect 11133 465 11171 499
rect 11205 465 11243 499
rect 11277 465 11315 499
rect 11349 465 11387 499
rect 11421 465 11459 499
rect 11493 465 11531 499
rect 11565 465 11603 499
rect 11637 465 11675 499
rect 11709 465 11747 499
rect 11781 465 11819 499
rect 11853 465 11891 499
rect 11925 465 11963 499
rect 11997 465 12035 499
rect 12069 465 12107 499
rect 12141 465 12179 499
rect 12213 465 12251 499
rect 12285 465 12323 499
rect 12357 465 12395 499
rect 12429 465 12467 499
rect 12501 465 12539 499
rect 12573 465 12611 499
rect 12645 465 12683 499
rect 12717 465 12755 499
rect 12789 465 12827 499
rect 12861 465 12899 499
rect 12933 465 12971 499
rect 13005 465 13043 499
rect 13077 465 13115 499
rect 13149 465 13187 499
rect 13221 465 13259 499
rect 13293 465 13331 499
rect 13365 465 13403 499
rect 13437 465 13475 499
rect 13509 465 13547 499
rect 13581 465 13619 499
rect 13653 465 13691 499
rect 13725 465 13763 499
rect 13797 465 13835 499
rect 13869 465 13907 499
rect 13941 465 13979 499
rect 14013 465 14051 499
rect 14085 465 14123 499
rect 14157 465 14195 499
rect 14229 465 14267 499
rect 14301 465 14339 499
rect 14373 465 14411 499
rect 14445 481 14483 499
rect 14517 481 14555 499
rect 14589 481 14627 499
rect 14661 481 14699 499
rect 14733 481 14771 499
rect 14445 465 14465 481
rect 14517 465 14539 481
rect 14589 465 14613 481
rect 14661 465 14686 481
rect 14733 465 14759 481
rect 14805 465 14843 499
rect 14877 465 14907 499
rect 229 463 343 465
rect 377 463 419 465
rect 453 463 495 465
rect 529 463 571 465
rect 605 463 648 465
rect 682 463 14465 465
rect 229 447 14465 463
rect 14499 447 14539 465
rect 14573 447 14613 465
rect 14647 447 14686 465
rect 14720 447 14759 465
rect 14793 447 14907 465
rect 229 431 14907 447
rect 229 397 302 431
rect 336 397 375 431
rect 409 397 448 431
rect 482 397 521 431
rect 555 397 594 431
rect 628 397 667 431
rect 701 397 740 431
rect 774 397 813 431
rect 847 397 886 431
rect 920 397 959 431
rect 993 397 1032 431
rect 1066 397 1105 431
rect 1139 397 1178 431
rect 1212 397 1251 431
rect 1285 397 1324 431
rect 1358 397 1397 431
rect 1431 397 1470 431
rect 1504 397 1543 431
rect 1577 397 1616 431
rect 1650 397 1689 431
rect 1723 397 1762 431
rect 1796 397 1835 431
rect 1869 397 1908 431
rect 1942 397 1981 431
rect 2015 397 2054 431
rect 2088 397 2127 431
rect 2161 397 2200 431
rect 2234 397 2273 431
rect 2307 397 2346 431
rect 2380 397 2419 431
rect 2453 397 2492 431
rect 2526 397 2565 431
rect 2599 397 2638 431
rect 2672 397 2711 431
rect 2745 397 2784 431
rect 2818 397 2857 431
rect 2891 397 2930 431
rect 2964 397 3003 431
rect 3037 397 3076 431
rect 3110 397 3149 431
rect 3183 397 3222 431
rect 3256 397 3295 431
rect 3329 397 3368 431
rect 3402 397 3441 431
rect 3475 397 3514 431
rect 3548 397 3587 431
rect 3621 397 3660 431
rect 3694 397 3733 431
rect 3767 397 3806 431
rect 3840 397 3879 431
rect 3913 397 3952 431
rect 3986 397 4025 431
rect 4059 397 4098 431
rect 4132 397 4171 431
rect 4205 397 4244 431
rect 4278 397 4317 431
rect 4351 397 4390 431
rect 4424 397 4463 431
rect 4497 397 4536 431
rect 4570 397 4609 431
rect 4643 397 4682 431
rect 4716 397 4755 431
rect 4789 397 4828 431
rect 4862 397 4901 431
rect 4935 397 4974 431
rect 5008 397 5047 431
rect 5081 397 5119 431
rect 5153 397 5191 431
rect 5225 397 5263 431
rect 5297 397 5335 431
rect 5369 397 5407 431
rect 5441 397 5479 431
rect 5513 397 5551 431
rect 5585 397 5623 431
rect 5657 397 5695 431
rect 5729 397 5767 431
rect 5801 397 5839 431
rect 5873 397 5911 431
rect 5945 397 5983 431
rect 6017 397 6055 431
rect 6089 397 6127 431
rect 6161 397 6199 431
rect 6233 397 6271 431
rect 6305 397 6343 431
rect 6377 397 6415 431
rect 6449 397 6487 431
rect 6521 397 6559 431
rect 6593 397 6631 431
rect 6665 397 6703 431
rect 6737 397 6775 431
rect 6809 397 6847 431
rect 6881 397 6919 431
rect 6953 397 6991 431
rect 7025 397 7063 431
rect 7097 397 7135 431
rect 7169 397 7207 431
rect 7241 397 7279 431
rect 7313 397 7351 431
rect 7385 397 7423 431
rect 7457 397 7495 431
rect 7529 397 7567 431
rect 7601 397 7639 431
rect 7673 397 7711 431
rect 7745 397 7783 431
rect 7817 397 7855 431
rect 7889 397 7927 431
rect 7961 397 7999 431
rect 8033 397 8071 431
rect 8105 397 8143 431
rect 8177 397 8215 431
rect 8249 397 8287 431
rect 8321 397 8359 431
rect 8393 397 8431 431
rect 8465 397 8503 431
rect 8537 397 8575 431
rect 8609 397 8647 431
rect 8681 397 8719 431
rect 8753 397 8791 431
rect 8825 397 8863 431
rect 8897 397 8935 431
rect 8969 397 9007 431
rect 9041 397 9079 431
rect 9113 397 9151 431
rect 9185 397 9223 431
rect 9257 397 9295 431
rect 9329 397 9367 431
rect 9401 397 9439 431
rect 9473 397 9511 431
rect 9545 397 9583 431
rect 9617 397 9655 431
rect 9689 397 9727 431
rect 9761 397 9799 431
rect 9833 397 9871 431
rect 9905 397 9943 431
rect 9977 397 10015 431
rect 10049 397 10087 431
rect 10121 397 10159 431
rect 10193 397 10231 431
rect 10265 397 10303 431
rect 10337 397 10375 431
rect 10409 397 10447 431
rect 10481 397 10519 431
rect 10553 397 10591 431
rect 10625 397 10663 431
rect 10697 397 10735 431
rect 10769 397 10807 431
rect 10841 397 10879 431
rect 10913 397 10951 431
rect 10985 397 11023 431
rect 11057 397 11095 431
rect 11129 397 11167 431
rect 11201 397 11239 431
rect 11273 397 11311 431
rect 11345 397 11383 431
rect 11417 397 11455 431
rect 11489 397 11527 431
rect 11561 397 11599 431
rect 11633 397 11671 431
rect 11705 397 11743 431
rect 11777 397 11815 431
rect 11849 397 11887 431
rect 11921 397 11959 431
rect 11993 397 12031 431
rect 12065 397 12103 431
rect 12137 397 12175 431
rect 12209 397 12247 431
rect 12281 397 12319 431
rect 12353 397 12391 431
rect 12425 397 12463 431
rect 12497 397 12535 431
rect 12569 397 12607 431
rect 12641 397 12679 431
rect 12713 397 12751 431
rect 12785 397 12823 431
rect 12857 397 12895 431
rect 12929 397 12967 431
rect 13001 397 13039 431
rect 13073 397 13111 431
rect 13145 397 13183 431
rect 13217 397 13255 431
rect 13289 397 13327 431
rect 13361 397 13399 431
rect 13433 397 13471 431
rect 13505 397 13543 431
rect 13577 397 13615 431
rect 13649 397 13687 431
rect 13721 397 13759 431
rect 13793 397 13831 431
rect 13865 397 13903 431
rect 13937 397 13975 431
rect 14009 397 14047 431
rect 14081 397 14119 431
rect 14153 397 14191 431
rect 14225 397 14263 431
rect 14297 397 14335 431
rect 14369 397 14407 431
rect 14441 397 14479 431
rect 14513 397 14551 431
rect 14585 397 14623 431
rect 14657 397 14695 431
rect 14729 397 14767 431
rect 14801 397 14839 431
rect 14873 397 14907 431
rect 229 375 14907 397
rect 229 363 361 375
rect 395 363 434 375
rect 468 363 507 375
rect 541 363 580 375
rect 614 363 653 375
rect 687 363 726 375
rect 760 363 799 375
rect 833 363 872 375
rect 906 363 945 375
rect 979 363 1018 375
rect 1052 363 1091 375
rect 1125 363 1164 375
rect 1198 363 1237 375
rect 1271 363 1310 375
rect 1344 363 1383 375
rect 1417 363 1456 375
rect 1490 363 1529 375
rect 1563 363 1602 375
rect 1636 363 1675 375
rect 1709 363 1748 375
rect 1782 363 1821 375
rect 1855 363 1894 375
rect 1928 363 1967 375
rect 2001 363 2040 375
rect 2074 363 2113 375
rect 2147 363 2186 375
rect 2220 363 2259 375
rect 2293 363 2332 375
rect 2366 363 2405 375
rect 2439 363 2478 375
rect 2512 363 2551 375
rect 2585 363 2624 375
rect 2658 363 2697 375
rect 2731 363 2770 375
rect 2804 363 2843 375
rect 2877 363 2916 375
rect 2950 363 2989 375
rect 3023 363 3062 375
rect 3096 363 3135 375
rect 3169 363 3208 375
rect 3242 363 3281 375
rect 3315 363 3354 375
rect 3388 363 3427 375
rect 3461 363 3500 375
rect 3534 363 3573 375
rect 3607 363 3646 375
rect 3680 363 3719 375
rect 3753 363 3792 375
rect 3826 363 3865 375
rect 3899 363 3938 375
rect 3972 363 4011 375
rect 4045 363 4084 375
rect 4118 363 4157 375
rect 4191 363 4229 375
rect 4263 363 4301 375
rect 4335 363 4373 375
rect 4407 363 4445 375
rect 4479 363 4517 375
rect 4551 363 4589 375
rect 4623 363 4661 375
rect 4695 363 4733 375
rect 4767 363 4805 375
rect 4839 363 4877 375
rect 4911 363 4949 375
rect 4983 363 5021 375
rect 5055 363 5093 375
rect 5127 363 5165 375
rect 5199 363 5237 375
rect 5271 363 5309 375
rect 5343 363 5381 375
rect 5415 363 5453 375
rect 5487 363 5525 375
rect 5559 363 5597 375
rect 5631 363 5669 375
rect 5703 363 5741 375
rect 5775 363 5813 375
rect 5847 363 5885 375
rect 5919 363 5957 375
rect 5991 363 6029 375
rect 6063 363 6101 375
rect 6135 363 6173 375
rect 6207 363 6245 375
rect 6279 363 6317 375
rect 6351 363 6389 375
rect 6423 363 6461 375
rect 6495 363 6533 375
rect 6567 363 6605 375
rect 6639 363 6677 375
rect 6711 363 6749 375
rect 6783 363 6821 375
rect 6855 363 6893 375
rect 6927 363 6965 375
rect 6999 363 7037 375
rect 7071 363 7109 375
rect 7143 363 7181 375
rect 7215 363 7253 375
rect 7287 363 7325 375
rect 7359 363 7397 375
rect 7431 363 7469 375
rect 7503 363 7541 375
rect 7575 363 7613 375
rect 7647 363 7685 375
rect 7719 363 7757 375
rect 7791 363 7829 375
rect 7863 363 7901 375
rect 7935 363 7973 375
rect 8007 363 8045 375
rect 8079 363 8117 375
rect 8151 363 8189 375
rect 8223 363 8261 375
rect 8295 363 8333 375
rect 8367 363 8405 375
rect 8439 363 8477 375
rect 8511 363 8549 375
rect 8583 363 8621 375
rect 8655 363 8693 375
rect 8727 363 8765 375
rect 8799 363 8837 375
rect 8871 363 8909 375
rect 8943 363 8981 375
rect 9015 363 9053 375
rect 9087 363 9125 375
rect 9159 363 9197 375
rect 9231 363 9269 375
rect 9303 363 9341 375
rect 9375 363 9413 375
rect 9447 363 9485 375
rect 9519 363 9557 375
rect 9591 363 9629 375
rect 9663 363 9701 375
rect 9735 363 9773 375
rect 9807 363 9845 375
rect 9879 363 9917 375
rect 9951 363 9989 375
rect 10023 363 10061 375
rect 10095 363 10133 375
rect 10167 363 10205 375
rect 10239 363 10277 375
rect 10311 363 10349 375
rect 10383 363 10421 375
rect 10455 363 10493 375
rect 10527 363 10565 375
rect 10599 363 10637 375
rect 10671 363 10709 375
rect 10743 363 10781 375
rect 10815 363 10853 375
rect 10887 363 10925 375
rect 10959 363 10997 375
rect 11031 363 11069 375
rect 11103 363 11141 375
rect 11175 363 11213 375
rect 11247 363 11285 375
rect 11319 363 11357 375
rect 11391 363 11429 375
rect 11463 363 11501 375
rect 11535 363 11573 375
rect 11607 363 11645 375
rect 11679 363 11717 375
rect 11751 363 11789 375
rect 11823 363 11861 375
rect 11895 363 11933 375
rect 11967 363 12005 375
rect 12039 363 12077 375
rect 12111 363 12149 375
rect 12183 363 12221 375
rect 12255 363 12293 375
rect 12327 363 12365 375
rect 12399 363 12437 375
rect 12471 363 12509 375
rect 12543 363 12581 375
rect 12615 363 12653 375
rect 12687 363 12725 375
rect 12759 363 12797 375
rect 12831 363 12869 375
rect 12903 363 12941 375
rect 12975 363 13013 375
rect 13047 363 13085 375
rect 13119 363 13157 375
rect 13191 363 13229 375
rect 13263 363 13301 375
rect 13335 363 13373 375
rect 13407 363 13445 375
rect 13479 363 13517 375
rect 13551 363 13589 375
rect 13623 363 13661 375
rect 13695 363 13733 375
rect 13767 363 13805 375
rect 13839 363 13877 375
rect 13911 363 13949 375
rect 13983 363 14021 375
rect 14055 363 14093 375
rect 14127 363 14165 375
rect 14199 363 14237 375
rect 14271 363 14309 375
rect 14343 363 14381 375
rect 14415 363 14453 375
rect 14487 363 14525 375
rect 14559 363 14597 375
rect 14631 363 14669 375
rect 14703 363 14741 375
rect 14775 363 14907 375
rect 229 331 302 363
rect 36 329 302 331
rect 336 341 361 363
rect 409 341 434 363
rect 482 341 507 363
rect 555 341 580 363
rect 628 341 653 363
rect 701 341 726 363
rect 774 341 799 363
rect 847 341 872 363
rect 920 341 945 363
rect 993 341 1018 363
rect 1066 341 1091 363
rect 1139 341 1164 363
rect 1212 341 1237 363
rect 1285 341 1310 363
rect 1358 341 1383 363
rect 1431 341 1456 363
rect 1504 341 1529 363
rect 1577 341 1602 363
rect 1650 341 1675 363
rect 1723 341 1748 363
rect 1796 341 1821 363
rect 1869 341 1894 363
rect 1942 341 1967 363
rect 2015 341 2040 363
rect 2088 341 2113 363
rect 2161 341 2186 363
rect 2234 341 2259 363
rect 2307 341 2332 363
rect 2380 341 2405 363
rect 2453 341 2478 363
rect 2526 341 2551 363
rect 2599 341 2624 363
rect 2672 341 2697 363
rect 2745 341 2770 363
rect 2818 341 2843 363
rect 2891 341 2916 363
rect 2964 341 2989 363
rect 3037 341 3062 363
rect 3110 341 3135 363
rect 3183 341 3208 363
rect 3256 341 3281 363
rect 3329 341 3354 363
rect 3402 341 3427 363
rect 3474 341 3500 363
rect 3546 341 3573 363
rect 3618 341 3646 363
rect 3690 341 3719 363
rect 3762 341 3792 363
rect 3834 341 3865 363
rect 3906 341 3938 363
rect 3978 341 4011 363
rect 4050 341 4084 363
rect 4122 341 4157 363
rect 4194 341 4229 363
rect 4266 341 4301 363
rect 4338 341 4373 363
rect 4410 341 4445 363
rect 4482 341 4517 363
rect 4554 341 4589 363
rect 4626 341 4661 363
rect 4698 341 4733 363
rect 4770 341 4805 363
rect 4842 341 4877 363
rect 4914 341 4949 363
rect 4986 341 5021 363
rect 5058 341 5093 363
rect 5130 341 5165 363
rect 5202 341 5237 363
rect 5274 341 5309 363
rect 5346 341 5381 363
rect 5418 341 5453 363
rect 5490 341 5525 363
rect 5562 341 5597 363
rect 5634 341 5669 363
rect 5706 341 5741 363
rect 5778 341 5813 363
rect 5850 341 5885 363
rect 5922 341 5957 363
rect 5994 341 6029 363
rect 6066 341 6101 363
rect 6138 341 6173 363
rect 6210 341 6245 363
rect 6282 341 6317 363
rect 6354 341 6389 363
rect 6426 341 6461 363
rect 6498 341 6533 363
rect 6570 341 6605 363
rect 6642 341 6677 363
rect 6714 341 6749 363
rect 6786 341 6821 363
rect 6858 341 6893 363
rect 6930 341 6965 363
rect 7002 341 7037 363
rect 7074 341 7109 363
rect 7146 341 7181 363
rect 7218 341 7253 363
rect 7290 341 7325 363
rect 7362 341 7397 363
rect 7434 341 7469 363
rect 7506 341 7541 363
rect 7578 341 7613 363
rect 7650 341 7685 363
rect 7722 341 7757 363
rect 7794 341 7829 363
rect 7866 341 7901 363
rect 7938 341 7973 363
rect 8010 341 8045 363
rect 8082 341 8117 363
rect 8154 341 8189 363
rect 8226 341 8261 363
rect 8298 341 8333 363
rect 8370 341 8405 363
rect 8442 341 8477 363
rect 8514 341 8549 363
rect 8586 341 8621 363
rect 8658 341 8693 363
rect 8730 341 8765 363
rect 8802 341 8837 363
rect 8874 341 8909 363
rect 8946 341 8981 363
rect 9018 341 9053 363
rect 9090 341 9125 363
rect 9162 341 9197 363
rect 9234 341 9269 363
rect 9306 341 9341 363
rect 9378 341 9413 363
rect 9450 341 9485 363
rect 9522 341 9557 363
rect 9594 341 9629 363
rect 9666 341 9701 363
rect 9738 341 9773 363
rect 9810 341 9845 363
rect 9882 341 9917 363
rect 9954 341 9989 363
rect 10026 341 10061 363
rect 10098 341 10133 363
rect 10170 341 10205 363
rect 10242 341 10277 363
rect 10314 341 10349 363
rect 10386 341 10421 363
rect 10458 341 10493 363
rect 10530 341 10565 363
rect 10602 341 10637 363
rect 10674 341 10709 363
rect 10746 341 10781 363
rect 10818 341 10853 363
rect 10890 341 10925 363
rect 10962 341 10997 363
rect 11034 341 11069 363
rect 11106 341 11141 363
rect 11178 341 11213 363
rect 11250 341 11285 363
rect 11322 341 11357 363
rect 11394 341 11429 363
rect 11466 341 11501 363
rect 11538 341 11573 363
rect 11610 341 11645 363
rect 11682 341 11717 363
rect 11754 341 11789 363
rect 11826 341 11861 363
rect 11898 341 11933 363
rect 11970 341 12005 363
rect 12042 341 12077 363
rect 12114 341 12149 363
rect 12186 341 12221 363
rect 12258 341 12293 363
rect 12330 341 12365 363
rect 12402 341 12437 363
rect 12474 341 12509 363
rect 12546 341 12581 363
rect 12618 341 12653 363
rect 12690 341 12725 363
rect 12762 341 12797 363
rect 12834 341 12869 363
rect 12906 341 12941 363
rect 12978 341 13013 363
rect 13050 341 13085 363
rect 13122 341 13157 363
rect 13194 341 13229 363
rect 13266 341 13301 363
rect 13338 341 13373 363
rect 13410 341 13445 363
rect 13482 341 13517 363
rect 13554 341 13589 363
rect 13626 341 13661 363
rect 13698 341 13733 363
rect 13770 341 13805 363
rect 13842 341 13877 363
rect 13914 341 13949 363
rect 13986 341 14021 363
rect 14058 341 14093 363
rect 14130 341 14165 363
rect 14202 341 14237 363
rect 14274 341 14309 363
rect 14346 341 14381 363
rect 14418 341 14453 363
rect 14490 341 14525 363
rect 14562 341 14597 363
rect 14634 341 14669 363
rect 14706 341 14741 363
rect 336 329 375 341
rect 409 329 448 341
rect 482 329 521 341
rect 555 329 594 341
rect 628 329 667 341
rect 701 329 740 341
rect 774 329 813 341
rect 847 329 886 341
rect 920 329 959 341
rect 993 329 1032 341
rect 1066 329 1105 341
rect 1139 329 1178 341
rect 1212 329 1251 341
rect 1285 329 1324 341
rect 1358 329 1397 341
rect 1431 329 1470 341
rect 1504 329 1543 341
rect 1577 329 1616 341
rect 1650 329 1689 341
rect 1723 329 1762 341
rect 1796 329 1835 341
rect 1869 329 1908 341
rect 1942 329 1981 341
rect 2015 329 2054 341
rect 2088 329 2127 341
rect 2161 329 2200 341
rect 2234 329 2273 341
rect 2307 329 2346 341
rect 2380 329 2419 341
rect 2453 329 2492 341
rect 2526 329 2565 341
rect 2599 329 2638 341
rect 2672 329 2711 341
rect 2745 329 2784 341
rect 2818 329 2857 341
rect 2891 329 2930 341
rect 2964 329 3003 341
rect 3037 329 3076 341
rect 3110 329 3149 341
rect 3183 329 3222 341
rect 3256 329 3295 341
rect 3329 329 3368 341
rect 3402 329 3440 341
rect 3474 329 3512 341
rect 3546 329 3584 341
rect 3618 329 3656 341
rect 3690 329 3728 341
rect 3762 329 3800 341
rect 3834 329 3872 341
rect 3906 329 3944 341
rect 3978 329 4016 341
rect 4050 329 4088 341
rect 4122 329 4160 341
rect 4194 329 4232 341
rect 4266 329 4304 341
rect 4338 329 4376 341
rect 4410 329 4448 341
rect 4482 329 4520 341
rect 4554 329 4592 341
rect 4626 329 4664 341
rect 4698 329 4736 341
rect 4770 329 4808 341
rect 4842 329 4880 341
rect 4914 329 4952 341
rect 4986 329 5024 341
rect 5058 329 5096 341
rect 5130 329 5168 341
rect 5202 329 5240 341
rect 5274 329 5312 341
rect 5346 329 5384 341
rect 5418 329 5456 341
rect 5490 329 5528 341
rect 5562 329 5600 341
rect 5634 329 5672 341
rect 5706 329 5744 341
rect 5778 329 5816 341
rect 5850 329 5888 341
rect 5922 329 5960 341
rect 5994 329 6032 341
rect 6066 329 6104 341
rect 6138 329 6176 341
rect 6210 329 6248 341
rect 6282 329 6320 341
rect 6354 329 6392 341
rect 6426 329 6464 341
rect 6498 329 6536 341
rect 6570 329 6608 341
rect 6642 329 6680 341
rect 6714 329 6752 341
rect 6786 329 6824 341
rect 6858 329 6896 341
rect 6930 329 6968 341
rect 7002 329 7040 341
rect 7074 329 7112 341
rect 7146 329 7184 341
rect 7218 329 7256 341
rect 7290 329 7328 341
rect 7362 329 7400 341
rect 7434 329 7472 341
rect 7506 329 7544 341
rect 7578 329 7616 341
rect 7650 329 7688 341
rect 7722 329 7760 341
rect 7794 329 7832 341
rect 7866 329 7904 341
rect 7938 329 7976 341
rect 8010 329 8048 341
rect 8082 329 8120 341
rect 8154 329 8192 341
rect 8226 329 8264 341
rect 8298 329 8336 341
rect 8370 329 8408 341
rect 8442 329 8480 341
rect 8514 329 8552 341
rect 8586 329 8624 341
rect 8658 329 8696 341
rect 8730 329 8768 341
rect 8802 329 8840 341
rect 8874 329 8912 341
rect 8946 329 8984 341
rect 9018 329 9056 341
rect 9090 329 9128 341
rect 9162 329 9200 341
rect 9234 329 9272 341
rect 9306 329 9344 341
rect 9378 329 9416 341
rect 9450 329 9488 341
rect 9522 329 9560 341
rect 9594 329 9632 341
rect 9666 329 9704 341
rect 9738 329 9776 341
rect 9810 329 9848 341
rect 9882 329 9920 341
rect 9954 329 9992 341
rect 10026 329 10064 341
rect 10098 329 10136 341
rect 10170 329 10208 341
rect 10242 329 10280 341
rect 10314 329 10352 341
rect 10386 329 10424 341
rect 10458 329 10496 341
rect 10530 329 10568 341
rect 10602 329 10640 341
rect 10674 329 10712 341
rect 10746 329 10784 341
rect 10818 329 10856 341
rect 10890 329 10928 341
rect 10962 329 11000 341
rect 11034 329 11072 341
rect 11106 329 11144 341
rect 11178 329 11216 341
rect 11250 329 11288 341
rect 11322 329 11360 341
rect 11394 329 11432 341
rect 11466 329 11504 341
rect 11538 329 11576 341
rect 11610 329 11648 341
rect 11682 329 11720 341
rect 11754 329 11792 341
rect 11826 329 11864 341
rect 11898 329 11936 341
rect 11970 329 12008 341
rect 12042 329 12080 341
rect 12114 329 12152 341
rect 12186 329 12224 341
rect 12258 329 12296 341
rect 12330 329 12368 341
rect 12402 329 12440 341
rect 12474 329 12512 341
rect 12546 329 12584 341
rect 12618 329 12656 341
rect 12690 329 12728 341
rect 12762 329 12800 341
rect 12834 329 12872 341
rect 12906 329 12944 341
rect 12978 329 13016 341
rect 13050 329 13088 341
rect 13122 329 13160 341
rect 13194 329 13232 341
rect 13266 329 13304 341
rect 13338 329 13376 341
rect 13410 329 13448 341
rect 13482 329 13520 341
rect 13554 329 13592 341
rect 13626 329 13664 341
rect 13698 329 13736 341
rect 13770 329 13808 341
rect 13842 329 13880 341
rect 13914 329 13952 341
rect 13986 329 14024 341
rect 14058 329 14096 341
rect 14130 329 14168 341
rect 14202 329 14240 341
rect 14274 329 14312 341
rect 14346 329 14384 341
rect 14418 329 14456 341
rect 14490 329 14528 341
rect 14562 329 14600 341
rect 14634 329 14672 341
rect 14706 329 14744 341
rect 14778 329 14816 363
rect 14850 329 14888 363
rect 15085 348 15100 5062
rect 14922 329 14960 348
rect 14994 329 15100 348
rect 36 314 15100 329
<< viali >>
rect 361 5077 395 5111
rect 434 5077 468 5111
rect 507 5077 541 5111
rect 580 5077 614 5111
rect 653 5077 687 5111
rect 726 5077 760 5111
rect 799 5077 833 5111
rect 872 5077 906 5111
rect 945 5077 979 5111
rect 1018 5077 1052 5111
rect 1091 5077 1125 5111
rect 1164 5077 1198 5111
rect 1237 5077 1271 5111
rect 1310 5077 1344 5111
rect 1383 5077 1417 5111
rect 1456 5077 1490 5111
rect 1529 5077 1563 5111
rect 1602 5077 1636 5111
rect 1675 5077 1709 5111
rect 1748 5077 1782 5111
rect 1821 5077 1855 5111
rect 1894 5077 1928 5111
rect 1967 5077 2001 5111
rect 2040 5077 2074 5111
rect 2113 5077 2147 5111
rect 2186 5077 2220 5111
rect 2259 5077 2293 5111
rect 2332 5077 2366 5111
rect 2405 5077 2439 5111
rect 2478 5077 2512 5111
rect 2551 5077 2585 5111
rect 2624 5077 2658 5111
rect 2697 5077 2731 5111
rect 2770 5077 2804 5111
rect 2843 5077 2877 5111
rect 2916 5077 2950 5111
rect 2989 5077 3023 5111
rect 3062 5077 3096 5111
rect 3135 5077 3169 5111
rect 3208 5077 3242 5111
rect 3281 5077 3315 5111
rect 3354 5077 3388 5111
rect 3427 5077 3461 5111
rect 3500 5077 3534 5111
rect 3573 5077 3607 5111
rect 3646 5077 3680 5111
rect 3719 5077 3753 5111
rect 3792 5077 3826 5111
rect 3865 5077 3899 5111
rect 3938 5077 3972 5111
rect 4011 5077 4045 5111
rect 4084 5077 4118 5111
rect 4157 5077 4191 5111
rect 4229 5077 4263 5111
rect 4301 5077 4335 5111
rect 4373 5077 4407 5111
rect 4445 5077 4479 5111
rect 4517 5077 4551 5111
rect 4589 5077 4623 5111
rect 4661 5077 4695 5111
rect 4733 5077 4767 5111
rect 4805 5077 4839 5111
rect 4877 5077 4911 5111
rect 4949 5077 4983 5111
rect 5021 5077 5055 5111
rect 5093 5077 5127 5111
rect 5165 5077 5199 5111
rect 5237 5077 5271 5111
rect 5309 5077 5343 5111
rect 5381 5077 5415 5111
rect 5453 5077 5487 5111
rect 5525 5077 5559 5111
rect 5597 5077 5631 5111
rect 5669 5077 5703 5111
rect 5741 5077 5775 5111
rect 5813 5077 5847 5111
rect 5885 5077 5919 5111
rect 5957 5077 5991 5111
rect 6029 5077 6063 5111
rect 6101 5077 6135 5111
rect 6173 5077 6207 5111
rect 6245 5077 6279 5111
rect 6317 5077 6351 5111
rect 6389 5077 6423 5111
rect 6461 5077 6495 5111
rect 6533 5077 6567 5111
rect 6605 5077 6639 5111
rect 6677 5077 6711 5111
rect 6749 5077 6783 5111
rect 6821 5077 6855 5111
rect 6893 5077 6927 5111
rect 6965 5077 6999 5111
rect 7037 5077 7071 5111
rect 7109 5077 7143 5111
rect 7181 5077 7215 5111
rect 7253 5077 7287 5111
rect 7325 5077 7359 5111
rect 7397 5077 7431 5111
rect 7469 5077 7503 5111
rect 7541 5077 7575 5111
rect 7613 5077 7647 5111
rect 7685 5077 7719 5111
rect 7757 5077 7791 5111
rect 7829 5077 7863 5111
rect 7901 5077 7935 5111
rect 7973 5077 8007 5111
rect 8045 5077 8079 5111
rect 8117 5077 8151 5111
rect 8189 5077 8223 5111
rect 8261 5077 8295 5111
rect 8333 5077 8367 5111
rect 8405 5077 8439 5111
rect 8477 5077 8511 5111
rect 8549 5077 8583 5111
rect 8621 5077 8655 5111
rect 8693 5077 8727 5111
rect 8765 5077 8799 5111
rect 8837 5077 8871 5111
rect 8909 5077 8943 5111
rect 8981 5077 9015 5111
rect 9053 5077 9087 5111
rect 9125 5077 9159 5111
rect 9197 5077 9231 5111
rect 9269 5077 9303 5111
rect 9341 5077 9375 5111
rect 9413 5077 9447 5111
rect 9485 5077 9519 5111
rect 9557 5077 9591 5111
rect 9629 5077 9663 5111
rect 9701 5077 9735 5111
rect 9773 5077 9807 5111
rect 9845 5077 9879 5111
rect 9917 5077 9951 5111
rect 9989 5077 10023 5111
rect 10061 5077 10095 5111
rect 10133 5077 10167 5111
rect 10205 5077 10239 5111
rect 10277 5077 10311 5111
rect 10349 5077 10383 5111
rect 10421 5077 10455 5111
rect 10493 5077 10527 5111
rect 10565 5077 10599 5111
rect 10637 5077 10671 5111
rect 10709 5077 10743 5111
rect 10781 5077 10815 5111
rect 10853 5077 10887 5111
rect 10925 5077 10959 5111
rect 10997 5077 11031 5111
rect 11069 5077 11103 5111
rect 11141 5077 11175 5111
rect 11213 5077 11247 5111
rect 11285 5077 11319 5111
rect 11357 5077 11391 5111
rect 11429 5077 11463 5111
rect 11501 5077 11535 5111
rect 11573 5077 11607 5111
rect 11645 5077 11679 5111
rect 11717 5077 11751 5111
rect 11789 5077 11823 5111
rect 11861 5077 11895 5111
rect 11933 5077 11967 5111
rect 12005 5077 12039 5111
rect 12077 5077 12111 5111
rect 12149 5077 12183 5111
rect 12221 5077 12255 5111
rect 12293 5077 12327 5111
rect 12365 5077 12399 5111
rect 12437 5077 12471 5111
rect 12509 5077 12543 5111
rect 12581 5077 12615 5111
rect 12653 5077 12687 5111
rect 12725 5077 12759 5111
rect 12797 5077 12831 5111
rect 12869 5077 12903 5111
rect 12941 5077 12975 5111
rect 13013 5077 13047 5111
rect 13085 5077 13119 5111
rect 13157 5077 13191 5111
rect 13229 5077 13263 5111
rect 13301 5077 13335 5111
rect 13373 5077 13407 5111
rect 13445 5077 13479 5111
rect 13517 5077 13551 5111
rect 13589 5077 13623 5111
rect 13661 5077 13695 5111
rect 13733 5077 13767 5111
rect 13805 5077 13839 5111
rect 13877 5077 13911 5111
rect 13949 5077 13983 5111
rect 14021 5077 14055 5111
rect 14093 5077 14127 5111
rect 14165 5077 14199 5111
rect 14237 5077 14271 5111
rect 14309 5077 14343 5111
rect 14381 5077 14415 5111
rect 14453 5077 14487 5111
rect 14525 5077 14559 5111
rect 14597 5077 14631 5111
rect 14669 5077 14703 5111
rect 14741 5077 14775 5111
rect 51 5015 85 5045
rect 85 5034 142 5045
rect 142 5034 176 5045
rect 176 5034 214 5045
rect 214 5034 229 5045
rect 361 5034 392 5035
rect 392 5034 395 5035
rect 434 5034 464 5035
rect 464 5034 468 5035
rect 507 5034 536 5035
rect 536 5034 541 5035
rect 580 5034 608 5035
rect 608 5034 614 5035
rect 653 5034 680 5035
rect 680 5034 687 5035
rect 726 5034 752 5035
rect 752 5034 760 5035
rect 799 5034 824 5035
rect 824 5034 833 5035
rect 872 5034 896 5035
rect 896 5034 906 5035
rect 945 5034 968 5035
rect 968 5034 979 5035
rect 1018 5034 1040 5035
rect 1040 5034 1052 5035
rect 1091 5034 1112 5035
rect 1112 5034 1125 5035
rect 1164 5034 1184 5035
rect 1184 5034 1198 5035
rect 1237 5034 1256 5035
rect 1256 5034 1271 5035
rect 1310 5034 1328 5035
rect 1328 5034 1344 5035
rect 1383 5034 1400 5035
rect 1400 5034 1417 5035
rect 1456 5034 1472 5035
rect 1472 5034 1490 5035
rect 1529 5034 1544 5035
rect 1544 5034 1563 5035
rect 1602 5034 1616 5035
rect 1616 5034 1636 5035
rect 1675 5034 1688 5035
rect 1688 5034 1709 5035
rect 1748 5034 1760 5035
rect 1760 5034 1782 5035
rect 1821 5034 1832 5035
rect 1832 5034 1855 5035
rect 1894 5034 1904 5035
rect 1904 5034 1928 5035
rect 1967 5034 1976 5035
rect 1976 5034 2001 5035
rect 2040 5034 2048 5035
rect 2048 5034 2074 5035
rect 2113 5034 2120 5035
rect 2120 5034 2147 5035
rect 2186 5034 2192 5035
rect 2192 5034 2220 5035
rect 2259 5034 2264 5035
rect 2264 5034 2293 5035
rect 2332 5034 2336 5035
rect 2336 5034 2366 5035
rect 2405 5034 2408 5035
rect 2408 5034 2439 5035
rect 2478 5034 2480 5035
rect 2480 5034 2512 5035
rect 2551 5034 2552 5035
rect 2552 5034 2585 5035
rect 85 5015 229 5034
rect 51 5000 229 5015
rect 269 5000 303 5029
rect 361 5001 395 5034
rect 434 5001 468 5034
rect 507 5001 541 5034
rect 580 5001 614 5034
rect 653 5001 687 5034
rect 726 5001 760 5034
rect 799 5001 833 5034
rect 872 5001 906 5034
rect 945 5001 979 5034
rect 1018 5001 1052 5034
rect 1091 5001 1125 5034
rect 1164 5001 1198 5034
rect 1237 5001 1271 5034
rect 1310 5001 1344 5034
rect 1383 5001 1417 5034
rect 1456 5001 1490 5034
rect 1529 5001 1563 5034
rect 1602 5001 1636 5034
rect 1675 5001 1709 5034
rect 1748 5001 1782 5034
rect 1821 5001 1855 5034
rect 1894 5001 1928 5034
rect 1967 5001 2001 5034
rect 2040 5001 2074 5034
rect 2113 5001 2147 5034
rect 2186 5001 2220 5034
rect 2259 5001 2293 5034
rect 2332 5001 2366 5034
rect 2405 5001 2439 5034
rect 2478 5001 2512 5034
rect 2551 5001 2585 5034
rect 2624 5001 2658 5035
rect 2697 5001 2731 5035
rect 2770 5001 2804 5035
rect 2843 5001 2877 5035
rect 2916 5001 2950 5035
rect 2989 5034 3022 5035
rect 3022 5034 3023 5035
rect 3062 5034 3094 5035
rect 3094 5034 3096 5035
rect 3135 5034 3166 5035
rect 3166 5034 3169 5035
rect 3208 5034 3238 5035
rect 3238 5034 3242 5035
rect 3281 5034 3310 5035
rect 3310 5034 3315 5035
rect 3354 5034 3382 5035
rect 3382 5034 3388 5035
rect 3427 5034 3454 5035
rect 3454 5034 3461 5035
rect 3500 5034 3526 5035
rect 3526 5034 3534 5035
rect 3573 5034 3598 5035
rect 3598 5034 3607 5035
rect 3646 5034 3670 5035
rect 3670 5034 3680 5035
rect 3719 5034 3742 5035
rect 3742 5034 3753 5035
rect 3792 5034 3814 5035
rect 3814 5034 3826 5035
rect 3865 5034 3886 5035
rect 3886 5034 3899 5035
rect 3938 5034 3958 5035
rect 3958 5034 3972 5035
rect 4011 5034 4030 5035
rect 4030 5034 4045 5035
rect 4084 5034 4102 5035
rect 4102 5034 4118 5035
rect 4157 5034 4174 5035
rect 4174 5034 4191 5035
rect 4229 5034 4246 5035
rect 4246 5034 4263 5035
rect 4301 5034 4318 5035
rect 4318 5034 4335 5035
rect 4373 5034 4390 5035
rect 4390 5034 4407 5035
rect 4445 5034 4462 5035
rect 4462 5034 4479 5035
rect 4517 5034 4534 5035
rect 4534 5034 4551 5035
rect 4589 5034 4606 5035
rect 4606 5034 4623 5035
rect 4661 5034 4678 5035
rect 4678 5034 4695 5035
rect 4733 5034 4750 5035
rect 4750 5034 4767 5035
rect 4805 5034 4822 5035
rect 4822 5034 4839 5035
rect 4877 5034 4894 5035
rect 4894 5034 4911 5035
rect 4949 5034 4966 5035
rect 4966 5034 4983 5035
rect 5021 5034 5038 5035
rect 5038 5034 5055 5035
rect 5093 5034 5110 5035
rect 5110 5034 5127 5035
rect 5165 5034 5182 5035
rect 5182 5034 5199 5035
rect 5237 5034 5254 5035
rect 5254 5034 5271 5035
rect 5309 5034 5326 5035
rect 5326 5034 5343 5035
rect 5381 5034 5398 5035
rect 5398 5034 5415 5035
rect 5453 5034 5470 5035
rect 5470 5034 5487 5035
rect 5525 5034 5542 5035
rect 5542 5034 5559 5035
rect 5597 5034 5614 5035
rect 5614 5034 5631 5035
rect 5669 5034 5686 5035
rect 5686 5034 5703 5035
rect 5741 5034 5758 5035
rect 5758 5034 5775 5035
rect 5813 5034 5830 5035
rect 5830 5034 5847 5035
rect 5885 5034 5902 5035
rect 5902 5034 5919 5035
rect 5957 5034 5974 5035
rect 5974 5034 5991 5035
rect 6029 5034 6046 5035
rect 6046 5034 6063 5035
rect 6101 5034 6118 5035
rect 6118 5034 6135 5035
rect 6173 5034 6190 5035
rect 6190 5034 6207 5035
rect 6245 5034 6262 5035
rect 6262 5034 6279 5035
rect 6317 5034 6334 5035
rect 6334 5034 6351 5035
rect 6389 5034 6406 5035
rect 6406 5034 6423 5035
rect 6461 5034 6478 5035
rect 6478 5034 6495 5035
rect 6533 5034 6550 5035
rect 6550 5034 6567 5035
rect 6605 5034 6622 5035
rect 6622 5034 6639 5035
rect 6677 5034 6694 5035
rect 6694 5034 6711 5035
rect 6749 5034 6766 5035
rect 6766 5034 6783 5035
rect 6821 5034 6838 5035
rect 6838 5034 6855 5035
rect 6893 5034 6910 5035
rect 6910 5034 6927 5035
rect 6965 5034 6982 5035
rect 6982 5034 6999 5035
rect 7037 5034 7054 5035
rect 7054 5034 7071 5035
rect 7109 5034 7126 5035
rect 7126 5034 7143 5035
rect 7181 5034 7198 5035
rect 7198 5034 7215 5035
rect 7253 5034 7270 5035
rect 7270 5034 7287 5035
rect 7325 5034 7342 5035
rect 7342 5034 7359 5035
rect 7397 5034 7414 5035
rect 7414 5034 7431 5035
rect 7469 5034 7486 5035
rect 7486 5034 7503 5035
rect 7541 5034 7558 5035
rect 7558 5034 7575 5035
rect 7613 5034 7630 5035
rect 7630 5034 7647 5035
rect 7685 5034 7702 5035
rect 7702 5034 7719 5035
rect 7757 5034 7774 5035
rect 7774 5034 7791 5035
rect 7829 5034 7846 5035
rect 7846 5034 7863 5035
rect 7901 5034 7918 5035
rect 7918 5034 7935 5035
rect 7973 5034 7990 5035
rect 7990 5034 8007 5035
rect 8045 5034 8062 5035
rect 8062 5034 8079 5035
rect 8117 5034 8134 5035
rect 8134 5034 8151 5035
rect 8189 5034 8206 5035
rect 8206 5034 8223 5035
rect 8261 5034 8278 5035
rect 8278 5034 8295 5035
rect 8333 5034 8350 5035
rect 8350 5034 8367 5035
rect 8405 5034 8422 5035
rect 8422 5034 8439 5035
rect 8477 5034 8494 5035
rect 8494 5034 8511 5035
rect 8549 5034 8566 5035
rect 8566 5034 8583 5035
rect 8621 5034 8638 5035
rect 8638 5034 8655 5035
rect 8693 5034 8710 5035
rect 8710 5034 8727 5035
rect 8765 5034 8782 5035
rect 8782 5034 8799 5035
rect 8837 5034 8854 5035
rect 8854 5034 8871 5035
rect 8909 5034 8926 5035
rect 8926 5034 8943 5035
rect 8981 5034 8998 5035
rect 8998 5034 9015 5035
rect 9053 5034 9070 5035
rect 9070 5034 9087 5035
rect 9125 5034 9142 5035
rect 9142 5034 9159 5035
rect 9197 5034 9214 5035
rect 9214 5034 9231 5035
rect 9269 5034 9286 5035
rect 9286 5034 9303 5035
rect 9341 5034 9358 5035
rect 9358 5034 9375 5035
rect 9413 5034 9430 5035
rect 9430 5034 9447 5035
rect 9485 5034 9502 5035
rect 9502 5034 9519 5035
rect 9557 5034 9574 5035
rect 9574 5034 9591 5035
rect 9629 5034 9646 5035
rect 9646 5034 9663 5035
rect 9701 5034 9718 5035
rect 9718 5034 9735 5035
rect 9773 5034 9790 5035
rect 9790 5034 9807 5035
rect 9845 5034 9862 5035
rect 9862 5034 9879 5035
rect 9917 5034 9934 5035
rect 9934 5034 9951 5035
rect 9989 5034 10006 5035
rect 10006 5034 10023 5035
rect 10061 5034 10078 5035
rect 10078 5034 10095 5035
rect 10133 5034 10151 5035
rect 10151 5034 10167 5035
rect 10205 5034 10224 5035
rect 10224 5034 10239 5035
rect 10277 5034 10297 5035
rect 10297 5034 10311 5035
rect 10349 5034 10370 5035
rect 10370 5034 10383 5035
rect 10421 5034 10443 5035
rect 10443 5034 10455 5035
rect 10493 5034 10516 5035
rect 10516 5034 10527 5035
rect 10565 5034 10589 5035
rect 10589 5034 10599 5035
rect 10637 5034 10662 5035
rect 10662 5034 10671 5035
rect 10709 5034 10735 5035
rect 10735 5034 10743 5035
rect 10781 5034 10808 5035
rect 10808 5034 10815 5035
rect 10853 5034 10881 5035
rect 10881 5034 10887 5035
rect 10925 5034 10954 5035
rect 10954 5034 10959 5035
rect 10997 5034 11027 5035
rect 11027 5034 11031 5035
rect 11069 5034 11100 5035
rect 11100 5034 11103 5035
rect 11141 5034 11173 5035
rect 11173 5034 11175 5035
rect 11213 5034 11246 5035
rect 11246 5034 11247 5035
rect 2989 5001 3023 5034
rect 3062 5001 3096 5034
rect 3135 5001 3169 5034
rect 3208 5001 3242 5034
rect 3281 5001 3315 5034
rect 3354 5001 3388 5034
rect 3427 5001 3461 5034
rect 3500 5001 3534 5034
rect 3573 5001 3607 5034
rect 3646 5001 3680 5034
rect 3719 5001 3753 5034
rect 3792 5001 3826 5034
rect 3865 5001 3899 5034
rect 3938 5001 3972 5034
rect 4011 5001 4045 5034
rect 4084 5001 4118 5034
rect 4157 5001 4191 5034
rect 4229 5001 4263 5034
rect 4301 5001 4335 5034
rect 4373 5001 4407 5034
rect 4445 5001 4479 5034
rect 4517 5001 4551 5034
rect 4589 5001 4623 5034
rect 4661 5001 4695 5034
rect 4733 5001 4767 5034
rect 4805 5001 4839 5034
rect 4877 5001 4911 5034
rect 4949 5001 4983 5034
rect 5021 5001 5055 5034
rect 5093 5001 5127 5034
rect 5165 5001 5199 5034
rect 5237 5001 5271 5034
rect 5309 5001 5343 5034
rect 5381 5001 5415 5034
rect 5453 5001 5487 5034
rect 5525 5001 5559 5034
rect 5597 5001 5631 5034
rect 5669 5001 5703 5034
rect 5741 5001 5775 5034
rect 5813 5001 5847 5034
rect 5885 5001 5919 5034
rect 5957 5001 5991 5034
rect 6029 5001 6063 5034
rect 6101 5001 6135 5034
rect 6173 5001 6207 5034
rect 6245 5001 6279 5034
rect 6317 5001 6351 5034
rect 6389 5001 6423 5034
rect 6461 5001 6495 5034
rect 6533 5001 6567 5034
rect 6605 5001 6639 5034
rect 6677 5001 6711 5034
rect 6749 5001 6783 5034
rect 6821 5001 6855 5034
rect 6893 5001 6927 5034
rect 6965 5001 6999 5034
rect 7037 5001 7071 5034
rect 7109 5001 7143 5034
rect 7181 5001 7215 5034
rect 7253 5001 7287 5034
rect 7325 5001 7359 5034
rect 7397 5001 7431 5034
rect 7469 5001 7503 5034
rect 7541 5001 7575 5034
rect 7613 5001 7647 5034
rect 7685 5001 7719 5034
rect 7757 5001 7791 5034
rect 7829 5001 7863 5034
rect 7901 5001 7935 5034
rect 7973 5001 8007 5034
rect 8045 5001 8079 5034
rect 8117 5001 8151 5034
rect 8189 5001 8223 5034
rect 8261 5001 8295 5034
rect 8333 5001 8367 5034
rect 8405 5001 8439 5034
rect 8477 5001 8511 5034
rect 8549 5001 8583 5034
rect 8621 5001 8655 5034
rect 8693 5001 8727 5034
rect 8765 5001 8799 5034
rect 8837 5001 8871 5034
rect 8909 5001 8943 5034
rect 8981 5001 9015 5034
rect 9053 5001 9087 5034
rect 9125 5001 9159 5034
rect 9197 5001 9231 5034
rect 9269 5001 9303 5034
rect 9341 5001 9375 5034
rect 9413 5001 9447 5034
rect 9485 5001 9519 5034
rect 9557 5001 9591 5034
rect 9629 5001 9663 5034
rect 9701 5001 9735 5034
rect 9773 5001 9807 5034
rect 9845 5001 9879 5034
rect 9917 5001 9951 5034
rect 9989 5001 10023 5034
rect 10061 5001 10095 5034
rect 10133 5001 10167 5034
rect 10205 5001 10239 5034
rect 10277 5001 10311 5034
rect 10349 5001 10383 5034
rect 10421 5001 10455 5034
rect 10493 5001 10527 5034
rect 10565 5001 10599 5034
rect 10637 5001 10671 5034
rect 10709 5001 10743 5034
rect 10781 5001 10815 5034
rect 10853 5001 10887 5034
rect 10925 5001 10959 5034
rect 10997 5001 11031 5034
rect 11069 5001 11103 5034
rect 11141 5001 11175 5034
rect 11213 5001 11247 5034
rect 11285 5001 11319 5035
rect 11357 5001 11391 5035
rect 11429 5001 11463 5035
rect 11501 5001 11535 5035
rect 11573 5001 11607 5035
rect 11645 5001 11679 5035
rect 11717 5034 11718 5035
rect 11718 5034 11751 5035
rect 11789 5034 11791 5035
rect 11791 5034 11823 5035
rect 11861 5034 11864 5035
rect 11864 5034 11895 5035
rect 11933 5034 11937 5035
rect 11937 5034 11967 5035
rect 12005 5034 12010 5035
rect 12010 5034 12039 5035
rect 12077 5034 12083 5035
rect 12083 5034 12111 5035
rect 12149 5034 12156 5035
rect 12156 5034 12183 5035
rect 12221 5034 12229 5035
rect 12229 5034 12255 5035
rect 12293 5034 12302 5035
rect 12302 5034 12327 5035
rect 12365 5034 12375 5035
rect 12375 5034 12399 5035
rect 12437 5034 12448 5035
rect 12448 5034 12471 5035
rect 12509 5034 12521 5035
rect 12521 5034 12543 5035
rect 12581 5034 12594 5035
rect 12594 5034 12615 5035
rect 12653 5034 12667 5035
rect 12667 5034 12687 5035
rect 12725 5034 12740 5035
rect 12740 5034 12759 5035
rect 12797 5034 12813 5035
rect 12813 5034 12831 5035
rect 12869 5034 12886 5035
rect 12886 5034 12903 5035
rect 12941 5034 12959 5035
rect 12959 5034 12975 5035
rect 13013 5034 13032 5035
rect 13032 5034 13047 5035
rect 13085 5034 13105 5035
rect 13105 5034 13119 5035
rect 13157 5034 13178 5035
rect 13178 5034 13191 5035
rect 13229 5034 13251 5035
rect 13251 5034 13263 5035
rect 13301 5034 13324 5035
rect 13324 5034 13335 5035
rect 13373 5034 13397 5035
rect 13397 5034 13407 5035
rect 13445 5034 13470 5035
rect 13470 5034 13479 5035
rect 13517 5034 13543 5035
rect 13543 5034 13551 5035
rect 13589 5034 13616 5035
rect 13616 5034 13623 5035
rect 13661 5034 13689 5035
rect 13689 5034 13695 5035
rect 13733 5034 13762 5035
rect 13762 5034 13767 5035
rect 13805 5034 13835 5035
rect 13835 5034 13839 5035
rect 13877 5034 13908 5035
rect 13908 5034 13911 5035
rect 13949 5034 13981 5035
rect 13981 5034 13983 5035
rect 14021 5034 14054 5035
rect 14054 5034 14055 5035
rect 11717 5001 11751 5034
rect 11789 5001 11823 5034
rect 11861 5001 11895 5034
rect 11933 5001 11967 5034
rect 12005 5001 12039 5034
rect 12077 5001 12111 5034
rect 12149 5001 12183 5034
rect 12221 5001 12255 5034
rect 12293 5001 12327 5034
rect 12365 5001 12399 5034
rect 12437 5001 12471 5034
rect 12509 5001 12543 5034
rect 12581 5001 12615 5034
rect 12653 5001 12687 5034
rect 12725 5001 12759 5034
rect 12797 5001 12831 5034
rect 12869 5001 12903 5034
rect 12941 5001 12975 5034
rect 13013 5001 13047 5034
rect 13085 5001 13119 5034
rect 13157 5001 13191 5034
rect 13229 5001 13263 5034
rect 13301 5001 13335 5034
rect 13373 5001 13407 5034
rect 13445 5001 13479 5034
rect 13517 5001 13551 5034
rect 13589 5001 13623 5034
rect 13661 5001 13695 5034
rect 13733 5001 13767 5034
rect 13805 5001 13839 5034
rect 13877 5001 13911 5034
rect 13949 5001 13983 5034
rect 14021 5001 14055 5034
rect 14093 5034 14127 5035
rect 14093 5001 14127 5034
rect 14165 5034 14166 5035
rect 14166 5034 14199 5035
rect 14237 5034 14239 5035
rect 14239 5034 14271 5035
rect 14309 5034 14312 5035
rect 14312 5034 14343 5035
rect 14381 5034 14385 5035
rect 14385 5034 14415 5035
rect 14453 5034 14458 5035
rect 14458 5034 14487 5035
rect 14525 5034 14531 5035
rect 14531 5034 14559 5035
rect 14597 5034 14604 5035
rect 14604 5034 14631 5035
rect 14669 5034 14677 5035
rect 14677 5034 14703 5035
rect 14741 5034 14750 5035
rect 14750 5034 14775 5035
rect 14165 5001 14199 5034
rect 14237 5001 14271 5034
rect 14309 5001 14343 5034
rect 14381 5001 14415 5034
rect 14453 5001 14487 5034
rect 14525 5001 14559 5034
rect 14597 5001 14631 5034
rect 14669 5001 14703 5034
rect 14741 5001 14775 5034
rect 14832 5000 14866 5030
rect 51 4976 119 5000
rect 51 4942 85 4976
rect 85 4966 119 4976
rect 119 4966 153 5000
rect 153 4966 191 5000
rect 191 4966 225 5000
rect 225 4966 229 5000
rect 269 4995 297 5000
rect 297 4995 303 5000
rect 14832 4996 14857 5000
rect 14857 4996 14866 5000
rect 14907 5017 15085 5062
rect 14907 4983 14915 5017
rect 14915 4983 14949 5017
rect 14949 4983 14983 5017
rect 14983 4983 15017 5017
rect 15017 4983 15051 5017
rect 15051 4983 15085 5017
rect 85 4942 229 4966
rect 51 4932 229 4942
rect 269 4932 303 4956
rect 361 4932 395 4959
rect 434 4932 468 4959
rect 507 4932 541 4959
rect 580 4932 614 4959
rect 51 4926 187 4932
rect 51 4903 119 4926
rect 51 4869 85 4903
rect 85 4892 119 4903
rect 119 4892 153 4926
rect 153 4898 187 4926
rect 187 4898 221 4932
rect 221 4898 229 4932
rect 269 4922 293 4932
rect 293 4922 303 4932
rect 361 4925 365 4932
rect 365 4925 395 4932
rect 434 4925 437 4932
rect 437 4925 468 4932
rect 507 4925 509 4932
rect 509 4925 541 4932
rect 580 4925 581 4932
rect 581 4925 614 4932
rect 653 4925 687 4959
rect 726 4925 760 4959
rect 799 4925 833 4959
rect 872 4925 906 4959
rect 945 4925 979 4959
rect 1018 4932 1052 4959
rect 1091 4932 1125 4959
rect 1164 4932 1198 4959
rect 1237 4932 1271 4959
rect 1310 4932 1344 4959
rect 1383 4932 1417 4959
rect 1456 4932 1490 4959
rect 1529 4932 1563 4959
rect 1602 4932 1636 4959
rect 1675 4932 1709 4959
rect 1748 4932 1782 4959
rect 1821 4932 1855 4959
rect 1894 4932 1928 4959
rect 1967 4932 2001 4959
rect 2040 4932 2074 4959
rect 2113 4932 2147 4959
rect 2186 4932 2220 4959
rect 2259 4932 2293 4959
rect 2332 4932 2366 4959
rect 2405 4932 2439 4959
rect 2478 4932 2512 4959
rect 2551 4932 2585 4959
rect 2624 4932 2658 4959
rect 2697 4932 2731 4959
rect 2770 4932 2804 4959
rect 2843 4932 2877 4959
rect 2916 4932 2950 4959
rect 2989 4932 3023 4959
rect 3062 4932 3096 4959
rect 3135 4932 3169 4959
rect 3208 4932 3242 4959
rect 3281 4932 3315 4959
rect 3354 4932 3388 4959
rect 3427 4932 3461 4959
rect 3500 4932 3534 4959
rect 3573 4932 3607 4959
rect 3646 4932 3680 4959
rect 3719 4932 3753 4959
rect 3792 4932 3826 4959
rect 3865 4932 3899 4959
rect 3938 4932 3972 4959
rect 4011 4932 4045 4959
rect 4084 4932 4118 4959
rect 4157 4932 4191 4959
rect 4229 4932 4263 4959
rect 4301 4932 4335 4959
rect 4373 4932 4407 4959
rect 4445 4932 4479 4959
rect 4517 4932 4551 4959
rect 4589 4932 4623 4959
rect 4661 4932 4695 4959
rect 4733 4932 4767 4959
rect 4805 4932 4839 4959
rect 4877 4932 4911 4959
rect 4949 4932 4983 4959
rect 5021 4932 5055 4959
rect 5093 4932 5127 4959
rect 5165 4932 5199 4959
rect 5237 4932 5271 4959
rect 5309 4932 5343 4959
rect 5381 4932 5415 4959
rect 5453 4932 5487 4959
rect 5525 4932 5559 4959
rect 5597 4932 5631 4959
rect 5669 4932 5703 4959
rect 5741 4932 5775 4959
rect 5813 4932 5847 4959
rect 5885 4932 5919 4959
rect 5957 4932 5991 4959
rect 6029 4932 6063 4959
rect 6101 4932 6135 4959
rect 6173 4932 6207 4959
rect 6245 4932 6279 4959
rect 6317 4932 6351 4959
rect 6389 4932 6423 4959
rect 6461 4932 6495 4959
rect 6533 4932 6567 4959
rect 6605 4932 6639 4959
rect 6677 4932 6711 4959
rect 6749 4932 6783 4959
rect 6821 4932 6855 4959
rect 6893 4932 6927 4959
rect 6965 4932 6999 4959
rect 7037 4932 7071 4959
rect 7109 4932 7143 4959
rect 7181 4932 7215 4959
rect 7253 4932 7287 4959
rect 7325 4932 7359 4959
rect 7397 4932 7431 4959
rect 7469 4932 7503 4959
rect 7541 4932 7575 4959
rect 7613 4932 7647 4959
rect 7685 4932 7719 4959
rect 7757 4932 7791 4959
rect 7829 4932 7863 4959
rect 7901 4932 7935 4959
rect 7973 4932 8007 4959
rect 8045 4932 8079 4959
rect 8117 4932 8151 4959
rect 8189 4932 8223 4959
rect 8261 4932 8295 4959
rect 8333 4932 8367 4959
rect 8405 4932 8439 4959
rect 8477 4932 8511 4959
rect 8549 4932 8583 4959
rect 8621 4932 8655 4959
rect 8693 4932 8727 4959
rect 8765 4932 8799 4959
rect 8837 4932 8871 4959
rect 8909 4932 8943 4959
rect 8981 4932 9015 4959
rect 9053 4932 9087 4959
rect 9125 4932 9159 4959
rect 9197 4932 9231 4959
rect 9269 4932 9303 4959
rect 9341 4932 9375 4959
rect 9413 4932 9447 4959
rect 9485 4932 9519 4959
rect 9557 4932 9591 4959
rect 9629 4932 9663 4959
rect 9701 4932 9735 4959
rect 9773 4932 9807 4959
rect 9845 4932 9879 4959
rect 9917 4932 9951 4959
rect 9989 4932 10023 4959
rect 10061 4932 10095 4959
rect 10133 4932 10167 4959
rect 10205 4932 10239 4959
rect 10277 4932 10311 4959
rect 10349 4932 10383 4959
rect 10421 4932 10455 4959
rect 10493 4932 10527 4959
rect 10565 4932 10599 4959
rect 10637 4932 10671 4959
rect 10709 4932 10743 4959
rect 10781 4932 10815 4959
rect 10853 4932 10887 4959
rect 10925 4932 10959 4959
rect 10997 4932 11031 4959
rect 11069 4932 11103 4959
rect 11141 4932 11175 4959
rect 11213 4932 11247 4959
rect 11285 4932 11319 4959
rect 11357 4932 11391 4959
rect 11429 4932 11463 4959
rect 11501 4932 11535 4959
rect 11573 4932 11607 4959
rect 11645 4932 11679 4959
rect 11717 4932 11751 4959
rect 11789 4932 11823 4959
rect 11861 4932 11895 4959
rect 11933 4932 11967 4959
rect 12005 4932 12039 4959
rect 12077 4932 12111 4959
rect 12149 4932 12183 4959
rect 12221 4932 12255 4959
rect 12293 4932 12327 4959
rect 12365 4932 12399 4959
rect 12437 4932 12471 4959
rect 12509 4932 12543 4959
rect 12581 4932 12615 4959
rect 12653 4932 12687 4959
rect 12725 4932 12759 4959
rect 12797 4932 12831 4959
rect 12869 4932 12903 4959
rect 12941 4932 12975 4959
rect 13013 4932 13047 4959
rect 13085 4932 13119 4959
rect 13157 4932 13191 4959
rect 13229 4932 13263 4959
rect 13301 4932 13335 4959
rect 13373 4932 13407 4959
rect 13445 4932 13479 4959
rect 13517 4932 13551 4959
rect 13589 4932 13623 4959
rect 13661 4932 13695 4959
rect 13733 4932 13767 4959
rect 13805 4932 13839 4959
rect 13877 4932 13911 4959
rect 13949 4932 13983 4959
rect 14021 4932 14055 4959
rect 1018 4925 1051 4932
rect 1051 4925 1052 4932
rect 1091 4925 1123 4932
rect 1123 4925 1125 4932
rect 1164 4925 1195 4932
rect 1195 4925 1198 4932
rect 1237 4925 1267 4932
rect 1267 4925 1271 4932
rect 1310 4925 1339 4932
rect 1339 4925 1344 4932
rect 1383 4925 1411 4932
rect 1411 4925 1417 4932
rect 1456 4925 1483 4932
rect 1483 4925 1490 4932
rect 1529 4925 1555 4932
rect 1555 4925 1563 4932
rect 1602 4925 1627 4932
rect 1627 4925 1636 4932
rect 1675 4925 1699 4932
rect 1699 4925 1709 4932
rect 1748 4925 1771 4932
rect 1771 4925 1782 4932
rect 1821 4925 1843 4932
rect 1843 4925 1855 4932
rect 1894 4925 1915 4932
rect 1915 4925 1928 4932
rect 1967 4925 1987 4932
rect 1987 4925 2001 4932
rect 2040 4925 2059 4932
rect 2059 4925 2074 4932
rect 2113 4925 2131 4932
rect 2131 4925 2147 4932
rect 2186 4925 2203 4932
rect 2203 4925 2220 4932
rect 2259 4925 2275 4932
rect 2275 4925 2293 4932
rect 2332 4925 2347 4932
rect 2347 4925 2366 4932
rect 2405 4925 2419 4932
rect 2419 4925 2439 4932
rect 2478 4925 2491 4932
rect 2491 4925 2512 4932
rect 2551 4925 2563 4932
rect 2563 4925 2585 4932
rect 2624 4925 2635 4932
rect 2635 4925 2658 4932
rect 2697 4925 2707 4932
rect 2707 4925 2731 4932
rect 2770 4925 2779 4932
rect 2779 4925 2804 4932
rect 2843 4925 2851 4932
rect 2851 4925 2877 4932
rect 2916 4925 2923 4932
rect 2923 4925 2950 4932
rect 2989 4925 2995 4932
rect 2995 4925 3023 4932
rect 3062 4925 3067 4932
rect 3067 4925 3096 4932
rect 3135 4925 3139 4932
rect 3139 4925 3169 4932
rect 3208 4925 3211 4932
rect 3211 4925 3242 4932
rect 3281 4925 3283 4932
rect 3283 4925 3315 4932
rect 3354 4925 3355 4932
rect 3355 4925 3388 4932
rect 3427 4925 3461 4932
rect 3500 4925 3533 4932
rect 3533 4925 3534 4932
rect 3573 4925 3605 4932
rect 3605 4925 3607 4932
rect 3646 4925 3677 4932
rect 3677 4925 3680 4932
rect 3719 4925 3749 4932
rect 3749 4925 3753 4932
rect 3792 4925 3821 4932
rect 3821 4925 3826 4932
rect 3865 4925 3893 4932
rect 3893 4925 3899 4932
rect 3938 4925 3965 4932
rect 3965 4925 3972 4932
rect 4011 4925 4037 4932
rect 4037 4925 4045 4932
rect 4084 4925 4109 4932
rect 4109 4925 4118 4932
rect 4157 4925 4181 4932
rect 4181 4925 4191 4932
rect 4229 4925 4253 4932
rect 4253 4925 4263 4932
rect 4301 4925 4325 4932
rect 4325 4925 4335 4932
rect 4373 4925 4397 4932
rect 4397 4925 4407 4932
rect 4445 4925 4469 4932
rect 4469 4925 4479 4932
rect 4517 4925 4541 4932
rect 4541 4925 4551 4932
rect 4589 4925 4613 4932
rect 4613 4925 4623 4932
rect 4661 4925 4685 4932
rect 4685 4925 4695 4932
rect 4733 4925 4757 4932
rect 4757 4925 4767 4932
rect 4805 4925 4829 4932
rect 4829 4925 4839 4932
rect 4877 4925 4901 4932
rect 4901 4925 4911 4932
rect 4949 4925 4973 4932
rect 4973 4925 4983 4932
rect 5021 4925 5045 4932
rect 5045 4925 5055 4932
rect 5093 4925 5117 4932
rect 5117 4925 5127 4932
rect 5165 4925 5189 4932
rect 5189 4925 5199 4932
rect 5237 4925 5261 4932
rect 5261 4925 5271 4932
rect 5309 4925 5333 4932
rect 5333 4925 5343 4932
rect 5381 4925 5405 4932
rect 5405 4925 5415 4932
rect 5453 4925 5477 4932
rect 5477 4925 5487 4932
rect 5525 4925 5549 4932
rect 5549 4925 5559 4932
rect 5597 4925 5621 4932
rect 5621 4925 5631 4932
rect 5669 4925 5693 4932
rect 5693 4925 5703 4932
rect 5741 4925 5765 4932
rect 5765 4925 5775 4932
rect 5813 4925 5837 4932
rect 5837 4925 5847 4932
rect 5885 4925 5909 4932
rect 5909 4925 5919 4932
rect 5957 4925 5981 4932
rect 5981 4925 5991 4932
rect 6029 4925 6053 4932
rect 6053 4925 6063 4932
rect 6101 4925 6125 4932
rect 6125 4925 6135 4932
rect 6173 4925 6197 4932
rect 6197 4925 6207 4932
rect 6245 4925 6269 4932
rect 6269 4925 6279 4932
rect 6317 4925 6341 4932
rect 6341 4925 6351 4932
rect 6389 4925 6413 4932
rect 6413 4925 6423 4932
rect 6461 4925 6485 4932
rect 6485 4925 6495 4932
rect 6533 4925 6557 4932
rect 6557 4925 6567 4932
rect 6605 4925 6629 4932
rect 6629 4925 6639 4932
rect 6677 4925 6701 4932
rect 6701 4925 6711 4932
rect 6749 4925 6773 4932
rect 6773 4925 6783 4932
rect 6821 4925 6845 4932
rect 6845 4925 6855 4932
rect 6893 4925 6917 4932
rect 6917 4925 6927 4932
rect 6965 4925 6989 4932
rect 6989 4925 6999 4932
rect 7037 4925 7061 4932
rect 7061 4925 7071 4932
rect 7109 4925 7133 4932
rect 7133 4925 7143 4932
rect 7181 4925 7205 4932
rect 7205 4925 7215 4932
rect 7253 4925 7277 4932
rect 7277 4925 7287 4932
rect 7325 4925 7349 4932
rect 7349 4925 7359 4932
rect 7397 4925 7421 4932
rect 7421 4925 7431 4932
rect 7469 4925 7493 4932
rect 7493 4925 7503 4932
rect 7541 4925 7565 4932
rect 7565 4925 7575 4932
rect 7613 4925 7637 4932
rect 7637 4925 7647 4932
rect 7685 4925 7709 4932
rect 7709 4925 7719 4932
rect 7757 4925 7781 4932
rect 7781 4925 7791 4932
rect 7829 4925 7853 4932
rect 7853 4925 7863 4932
rect 7901 4925 7925 4932
rect 7925 4925 7935 4932
rect 7973 4925 7997 4932
rect 7997 4925 8007 4932
rect 8045 4925 8069 4932
rect 8069 4925 8079 4932
rect 8117 4925 8141 4932
rect 8141 4925 8151 4932
rect 8189 4925 8213 4932
rect 8213 4925 8223 4932
rect 8261 4925 8285 4932
rect 8285 4925 8295 4932
rect 8333 4925 8357 4932
rect 8357 4925 8367 4932
rect 8405 4925 8429 4932
rect 8429 4925 8439 4932
rect 8477 4925 8501 4932
rect 8501 4925 8511 4932
rect 8549 4925 8573 4932
rect 8573 4925 8583 4932
rect 8621 4925 8645 4932
rect 8645 4925 8655 4932
rect 8693 4925 8717 4932
rect 8717 4925 8727 4932
rect 8765 4925 8789 4932
rect 8789 4925 8799 4932
rect 8837 4925 8861 4932
rect 8861 4925 8871 4932
rect 8909 4925 8933 4932
rect 8933 4925 8943 4932
rect 8981 4925 9005 4932
rect 9005 4925 9015 4932
rect 9053 4925 9077 4932
rect 9077 4925 9087 4932
rect 9125 4925 9149 4932
rect 9149 4925 9159 4932
rect 9197 4925 9221 4932
rect 9221 4925 9231 4932
rect 9269 4925 9293 4932
rect 9293 4925 9303 4932
rect 9341 4925 9365 4932
rect 9365 4925 9375 4932
rect 9413 4925 9437 4932
rect 9437 4925 9447 4932
rect 9485 4925 9509 4932
rect 9509 4925 9519 4932
rect 9557 4925 9581 4932
rect 9581 4925 9591 4932
rect 9629 4925 9653 4932
rect 9653 4925 9663 4932
rect 9701 4925 9725 4932
rect 9725 4925 9735 4932
rect 9773 4925 9797 4932
rect 9797 4925 9807 4932
rect 9845 4925 9869 4932
rect 9869 4925 9879 4932
rect 9917 4925 9941 4932
rect 9941 4925 9951 4932
rect 9989 4925 10013 4932
rect 10013 4925 10023 4932
rect 10061 4925 10085 4932
rect 10085 4925 10095 4932
rect 10133 4925 10157 4932
rect 10157 4925 10167 4932
rect 10205 4925 10229 4932
rect 10229 4925 10239 4932
rect 10277 4925 10301 4932
rect 10301 4925 10311 4932
rect 10349 4925 10373 4932
rect 10373 4925 10383 4932
rect 10421 4925 10445 4932
rect 10445 4925 10455 4932
rect 10493 4925 10517 4932
rect 10517 4925 10527 4932
rect 10565 4925 10589 4932
rect 10589 4925 10599 4932
rect 10637 4925 10661 4932
rect 10661 4925 10671 4932
rect 10709 4925 10733 4932
rect 10733 4925 10743 4932
rect 10781 4925 10805 4932
rect 10805 4925 10815 4932
rect 10853 4925 10877 4932
rect 10877 4925 10887 4932
rect 10925 4925 10949 4932
rect 10949 4925 10959 4932
rect 10997 4925 11021 4932
rect 11021 4925 11031 4932
rect 11069 4925 11093 4932
rect 11093 4925 11103 4932
rect 11141 4925 11165 4932
rect 11165 4925 11175 4932
rect 11213 4925 11237 4932
rect 11237 4925 11247 4932
rect 11285 4925 11309 4932
rect 11309 4925 11319 4932
rect 11357 4925 11381 4932
rect 11381 4925 11391 4932
rect 11429 4925 11453 4932
rect 11453 4925 11463 4932
rect 11501 4925 11525 4932
rect 11525 4925 11535 4932
rect 11573 4925 11597 4932
rect 11597 4925 11607 4932
rect 11645 4925 11669 4932
rect 11669 4925 11679 4932
rect 11717 4925 11741 4932
rect 11741 4925 11751 4932
rect 11789 4925 11813 4932
rect 11813 4925 11823 4932
rect 11861 4925 11885 4932
rect 11885 4925 11895 4932
rect 11933 4925 11957 4932
rect 11957 4925 11967 4932
rect 12005 4925 12029 4932
rect 12029 4925 12039 4932
rect 12077 4925 12101 4932
rect 12101 4925 12111 4932
rect 12149 4925 12173 4932
rect 12173 4925 12183 4932
rect 12221 4925 12245 4932
rect 12245 4925 12255 4932
rect 12293 4925 12317 4932
rect 12317 4925 12327 4932
rect 12365 4925 12389 4932
rect 12389 4925 12399 4932
rect 12437 4925 12461 4932
rect 12461 4925 12471 4932
rect 12509 4925 12533 4932
rect 12533 4925 12543 4932
rect 12581 4925 12605 4932
rect 12605 4925 12615 4932
rect 12653 4925 12677 4932
rect 12677 4925 12687 4932
rect 12725 4925 12749 4932
rect 12749 4925 12759 4932
rect 12797 4925 12821 4932
rect 12821 4925 12831 4932
rect 12869 4925 12893 4932
rect 12893 4925 12903 4932
rect 12941 4925 12965 4932
rect 12965 4925 12975 4932
rect 13013 4925 13037 4932
rect 13037 4925 13047 4932
rect 13085 4925 13109 4932
rect 13109 4925 13119 4932
rect 13157 4925 13181 4932
rect 13181 4925 13191 4932
rect 13229 4925 13253 4932
rect 13253 4925 13263 4932
rect 13301 4925 13325 4932
rect 13325 4925 13335 4932
rect 13373 4925 13397 4932
rect 13397 4925 13407 4932
rect 13445 4925 13470 4932
rect 13470 4925 13479 4932
rect 13517 4925 13543 4932
rect 13543 4925 13551 4932
rect 13589 4925 13616 4932
rect 13616 4925 13623 4932
rect 13661 4925 13689 4932
rect 13689 4925 13695 4932
rect 13733 4925 13762 4932
rect 13762 4925 13767 4932
rect 13805 4925 13835 4932
rect 13835 4925 13839 4932
rect 13877 4925 13908 4932
rect 13908 4925 13911 4932
rect 13949 4925 13981 4932
rect 13981 4925 13983 4932
rect 14021 4925 14054 4932
rect 14054 4925 14055 4932
rect 14093 4932 14127 4959
rect 14093 4925 14127 4932
rect 14165 4932 14199 4959
rect 14237 4932 14271 4959
rect 14309 4932 14343 4959
rect 14381 4932 14415 4959
rect 14453 4932 14487 4959
rect 14525 4932 14559 4959
rect 14597 4932 14631 4959
rect 14669 4932 14703 4959
rect 14741 4932 14775 4959
rect 14832 4932 14866 4958
rect 14165 4925 14166 4932
rect 14166 4925 14199 4932
rect 14237 4925 14239 4932
rect 14239 4925 14271 4932
rect 14309 4925 14312 4932
rect 14312 4925 14343 4932
rect 14381 4925 14385 4932
rect 14385 4925 14415 4932
rect 14453 4925 14458 4932
rect 14458 4925 14487 4932
rect 14525 4925 14531 4932
rect 14531 4925 14559 4932
rect 14597 4925 14604 4932
rect 14604 4925 14631 4932
rect 14669 4925 14677 4932
rect 14677 4925 14703 4932
rect 14741 4925 14750 4932
rect 14750 4925 14775 4932
rect 14832 4924 14857 4932
rect 14857 4924 14866 4932
rect 14907 4945 15085 4983
rect 14907 4911 14915 4945
rect 14915 4911 14949 4945
rect 14949 4911 14983 4945
rect 14983 4911 15017 4945
rect 15017 4911 15051 4945
rect 15051 4911 15085 4945
rect 153 4892 229 4898
rect 85 4869 229 4892
rect 51 4857 229 4869
rect 269 4859 303 4883
rect 51 4852 187 4857
rect 51 4830 119 4852
rect 51 4796 85 4830
rect 85 4818 119 4830
rect 119 4818 153 4852
rect 153 4823 187 4852
rect 187 4823 221 4857
rect 221 4823 229 4857
rect 269 4849 296 4859
rect 296 4849 303 4859
rect 153 4818 229 4823
rect 85 4796 229 4818
rect 51 4782 229 4796
rect 269 4791 303 4810
rect 51 4778 187 4782
rect 51 4757 119 4778
rect 51 4723 85 4757
rect 85 4744 119 4757
rect 119 4744 153 4778
rect 153 4748 187 4778
rect 187 4748 221 4782
rect 221 4748 229 4782
rect 269 4776 296 4791
rect 296 4776 303 4791
rect 153 4744 229 4748
rect 85 4723 229 4744
rect 269 4723 303 4737
rect 51 4707 229 4723
rect 51 4704 187 4707
rect 51 4684 119 4704
rect 51 4650 85 4684
rect 85 4670 119 4684
rect 119 4670 153 4704
rect 153 4673 187 4704
rect 187 4673 221 4707
rect 221 4673 229 4707
rect 269 4703 296 4723
rect 296 4703 303 4723
rect 153 4670 229 4673
rect 85 4650 229 4670
rect 269 4655 303 4664
rect 51 4632 229 4650
rect 51 4630 187 4632
rect 51 4611 119 4630
rect 51 4577 85 4611
rect 85 4596 119 4611
rect 119 4596 153 4630
rect 153 4598 187 4630
rect 187 4598 221 4632
rect 221 4598 229 4632
rect 269 4630 296 4655
rect 296 4630 303 4655
rect 14832 4859 14866 4886
rect 14907 4873 15085 4911
rect 14832 4852 14840 4859
rect 14840 4852 14866 4859
rect 14907 4839 14915 4873
rect 14915 4839 14949 4873
rect 14949 4839 14983 4873
rect 14983 4839 15017 4873
rect 15017 4839 15051 4873
rect 15051 4839 15085 4873
rect 14832 4791 14866 4814
rect 14907 4801 15085 4839
rect 14832 4780 14840 4791
rect 14840 4780 14866 4791
rect 14907 4767 14915 4801
rect 14915 4767 14949 4801
rect 14949 4767 14983 4801
rect 14983 4767 15017 4801
rect 15017 4767 15051 4801
rect 15051 4767 15085 4801
rect 14832 4723 14866 4742
rect 14907 4729 15085 4767
rect 14832 4708 14840 4723
rect 14840 4708 14866 4723
rect 14907 4695 14915 4729
rect 14915 4695 14949 4729
rect 14949 4695 14983 4729
rect 14983 4695 15017 4729
rect 15017 4695 15051 4729
rect 15051 4695 15085 4729
rect 153 4596 229 4598
rect 85 4577 229 4596
rect 269 4587 303 4591
rect 51 4557 229 4577
rect 51 4556 187 4557
rect 51 4538 119 4556
rect 51 4504 85 4538
rect 85 4522 119 4538
rect 119 4522 153 4556
rect 153 4523 187 4556
rect 187 4523 221 4557
rect 221 4523 229 4557
rect 269 4557 296 4587
rect 296 4557 303 4587
rect 153 4522 229 4523
rect 85 4504 229 4522
rect 51 4483 229 4504
rect 269 4485 296 4518
rect 296 4485 303 4518
rect 269 4484 303 4485
rect 51 4482 187 4483
rect 51 4465 119 4482
rect 51 4431 85 4465
rect 85 4448 119 4465
rect 119 4448 153 4482
rect 153 4449 187 4482
rect 187 4449 221 4483
rect 221 4449 229 4483
rect 153 4448 229 4449
rect 85 4431 229 4448
rect 51 4409 229 4431
rect 269 4417 296 4445
rect 296 4417 303 4445
rect 269 4411 303 4417
rect 51 4408 187 4409
rect 51 4393 119 4408
rect 51 4359 85 4393
rect 85 4374 119 4393
rect 119 4374 153 4408
rect 153 4375 187 4408
rect 187 4375 221 4409
rect 221 4375 229 4409
rect 153 4374 229 4375
rect 85 4359 229 4374
rect 51 4335 229 4359
rect 269 4349 296 4372
rect 296 4349 303 4372
rect 269 4338 303 4349
rect 51 4334 187 4335
rect 51 4321 119 4334
rect 51 4287 85 4321
rect 85 4300 119 4321
rect 119 4300 153 4334
rect 153 4301 187 4334
rect 187 4301 221 4335
rect 221 4301 229 4335
rect 153 4300 229 4301
rect 85 4287 229 4300
rect 51 4261 229 4287
rect 269 4281 296 4299
rect 296 4281 303 4299
rect 269 4265 303 4281
rect 51 4260 187 4261
rect 51 4249 119 4260
rect 51 4215 85 4249
rect 85 4226 119 4249
rect 119 4226 153 4260
rect 153 4227 187 4260
rect 187 4227 221 4261
rect 221 4227 229 4261
rect 153 4226 229 4227
rect 85 4215 229 4226
rect 51 4187 229 4215
rect 269 4213 296 4226
rect 296 4213 303 4226
rect 269 4192 303 4213
rect 51 4186 187 4187
rect 51 4177 119 4186
rect 51 4143 85 4177
rect 85 4152 119 4177
rect 119 4152 153 4186
rect 153 4153 187 4186
rect 187 4153 221 4187
rect 221 4153 229 4187
rect 153 4152 229 4153
rect 85 4143 229 4152
rect 269 4145 296 4153
rect 296 4145 303 4153
rect 51 4113 229 4143
rect 269 4119 303 4145
rect 51 4112 187 4113
rect 51 4105 119 4112
rect 51 4071 85 4105
rect 85 4078 119 4105
rect 119 4078 153 4112
rect 153 4079 187 4112
rect 187 4079 221 4113
rect 221 4079 229 4113
rect 153 4078 229 4079
rect 85 4071 229 4078
rect 269 4077 296 4080
rect 296 4077 303 4080
rect 51 4039 229 4071
rect 269 4046 303 4077
rect 51 4038 187 4039
rect 51 4033 119 4038
rect 51 3999 85 4033
rect 85 4004 119 4033
rect 119 4004 153 4038
rect 153 4005 187 4038
rect 187 4005 221 4039
rect 221 4005 229 4039
rect 153 4004 229 4005
rect 85 3999 229 4004
rect 51 3965 229 3999
rect 269 3975 303 4007
rect 51 3964 187 3965
rect 51 3961 119 3964
rect 51 3927 85 3961
rect 85 3930 119 3961
rect 119 3930 153 3964
rect 153 3931 187 3964
rect 187 3931 221 3965
rect 221 3931 229 3965
rect 269 3973 296 3975
rect 296 3973 303 3975
rect 153 3930 229 3931
rect 85 3927 229 3930
rect 51 3891 229 3927
rect 269 3907 303 3934
rect 51 3890 187 3891
rect 51 3889 119 3890
rect 51 3855 85 3889
rect 85 3856 119 3889
rect 119 3856 153 3890
rect 153 3857 187 3890
rect 187 3857 221 3891
rect 221 3857 229 3891
rect 269 3900 296 3907
rect 296 3900 303 3907
rect 153 3856 229 3857
rect 85 3855 229 3856
rect 51 3817 229 3855
rect 269 3839 303 3861
rect 51 3783 85 3817
rect 85 3783 119 3817
rect 119 3783 153 3817
rect 153 3783 187 3817
rect 187 3783 221 3817
rect 221 3783 229 3817
rect 269 3827 296 3839
rect 296 3827 303 3839
rect 51 3707 229 3783
rect 269 3771 303 3788
rect 269 3754 296 3771
rect 296 3754 303 3771
rect 51 3673 85 3707
rect 85 3673 119 3707
rect 119 3673 153 3707
rect 153 3673 187 3707
rect 187 3673 221 3707
rect 221 3673 229 3707
rect 269 3703 303 3715
rect 51 3634 229 3673
rect 269 3681 296 3703
rect 296 3681 303 3703
rect 269 3635 303 3642
rect 51 3600 85 3634
rect 85 3600 119 3634
rect 119 3600 153 3634
rect 153 3600 187 3634
rect 187 3600 221 3634
rect 221 3600 229 3634
rect 269 3608 296 3635
rect 296 3608 303 3635
rect 51 3562 229 3600
rect 269 3567 303 3569
rect 51 3528 85 3562
rect 85 3528 119 3562
rect 119 3528 153 3562
rect 153 3528 187 3562
rect 187 3528 221 3562
rect 221 3528 229 3562
rect 269 3535 296 3567
rect 296 3535 303 3567
rect 51 3490 229 3528
rect 51 3456 85 3490
rect 85 3456 119 3490
rect 119 3456 153 3490
rect 153 3456 187 3490
rect 187 3456 221 3490
rect 221 3456 229 3490
rect 269 3465 296 3496
rect 296 3465 303 3496
rect 269 3462 303 3465
rect 51 3418 229 3456
rect 51 3384 85 3418
rect 85 3384 119 3418
rect 119 3384 153 3418
rect 153 3384 187 3418
rect 187 3384 221 3418
rect 221 3384 229 3418
rect 269 3397 296 3423
rect 296 3397 303 3423
rect 269 3389 303 3397
rect 51 3346 229 3384
rect 51 3312 85 3346
rect 85 3312 119 3346
rect 119 3312 153 3346
rect 153 3312 187 3346
rect 187 3312 221 3346
rect 221 3312 229 3346
rect 269 3329 296 3350
rect 296 3329 303 3350
rect 269 3316 303 3329
rect 51 3274 229 3312
rect 51 3240 85 3274
rect 85 3240 119 3274
rect 119 3240 153 3274
rect 153 3240 187 3274
rect 187 3240 221 3274
rect 221 3240 229 3274
rect 269 3261 296 3277
rect 296 3261 303 3277
rect 269 3243 303 3261
rect 51 3202 229 3240
rect 51 3168 85 3202
rect 85 3168 119 3202
rect 119 3168 153 3202
rect 153 3168 187 3202
rect 187 3168 221 3202
rect 221 3168 229 3202
rect 269 3193 296 3204
rect 296 3193 303 3204
rect 269 3170 303 3193
rect 51 3130 229 3168
rect 51 3096 85 3130
rect 85 3096 119 3130
rect 119 3096 153 3130
rect 153 3096 187 3130
rect 187 3096 221 3130
rect 221 3096 229 3130
rect 269 3125 296 3131
rect 296 3125 303 3131
rect 269 3097 303 3125
rect 51 3058 229 3096
rect 51 3024 85 3058
rect 85 3024 119 3058
rect 119 3024 153 3058
rect 153 3024 187 3058
rect 187 3024 221 3058
rect 221 3024 229 3058
rect 269 3057 296 3058
rect 296 3057 303 3058
rect 269 3024 303 3057
rect 51 2986 229 3024
rect 51 2952 85 2986
rect 85 2952 119 2986
rect 119 2952 153 2986
rect 153 2952 187 2986
rect 187 2952 221 2986
rect 221 2952 229 2986
rect 269 2955 303 2985
rect 51 2914 229 2952
rect 269 2951 296 2955
rect 296 2951 303 2955
rect 51 2880 85 2914
rect 85 2880 119 2914
rect 119 2880 153 2914
rect 153 2880 187 2914
rect 187 2880 221 2914
rect 221 2880 229 2914
rect 269 2887 303 2912
rect 51 2842 229 2880
rect 269 2878 296 2887
rect 296 2878 303 2887
rect 51 2808 85 2842
rect 85 2808 119 2842
rect 119 2808 153 2842
rect 153 2808 187 2842
rect 187 2808 221 2842
rect 221 2808 229 2842
rect 269 2819 303 2839
rect 51 2770 229 2808
rect 269 2805 296 2819
rect 296 2805 303 2819
rect 51 2736 85 2770
rect 85 2736 119 2770
rect 119 2736 153 2770
rect 153 2736 187 2770
rect 187 2736 221 2770
rect 221 2736 229 2770
rect 269 2751 303 2766
rect 51 2698 229 2736
rect 269 2732 296 2751
rect 296 2732 303 2751
rect 51 2664 85 2698
rect 85 2664 119 2698
rect 119 2664 153 2698
rect 153 2664 187 2698
rect 187 2664 221 2698
rect 221 2664 229 2698
rect 269 2683 303 2693
rect 51 2626 229 2664
rect 269 2659 296 2683
rect 296 2659 303 2683
rect 51 2592 85 2626
rect 85 2592 119 2626
rect 119 2592 153 2626
rect 153 2592 187 2626
rect 187 2592 221 2626
rect 221 2592 229 2626
rect 269 2615 303 2620
rect 51 2554 229 2592
rect 269 2586 296 2615
rect 296 2586 303 2615
rect 51 2520 85 2554
rect 85 2520 119 2554
rect 119 2520 153 2554
rect 153 2520 187 2554
rect 187 2520 221 2554
rect 221 2520 229 2554
rect 51 2482 229 2520
rect 269 2513 296 2547
rect 296 2513 303 2547
rect 51 2448 85 2482
rect 85 2448 119 2482
rect 119 2448 153 2482
rect 153 2448 187 2482
rect 187 2448 221 2482
rect 221 2448 229 2482
rect 51 2410 229 2448
rect 269 2445 296 2474
rect 296 2445 303 2474
rect 269 2440 303 2445
rect 51 2376 85 2410
rect 85 2376 119 2410
rect 119 2376 153 2410
rect 153 2376 187 2410
rect 187 2376 221 2410
rect 221 2376 229 2410
rect 269 2377 296 2401
rect 296 2377 303 2401
rect 51 2338 229 2376
rect 269 2367 303 2377
rect 51 2304 85 2338
rect 85 2304 119 2338
rect 119 2304 153 2338
rect 153 2304 187 2338
rect 187 2304 221 2338
rect 221 2304 229 2338
rect 269 2309 296 2328
rect 296 2309 303 2328
rect 51 2266 229 2304
rect 269 2294 303 2309
rect 51 2232 85 2266
rect 85 2232 119 2266
rect 119 2232 153 2266
rect 153 2232 187 2266
rect 187 2232 221 2266
rect 221 2232 229 2266
rect 269 2241 296 2255
rect 296 2241 303 2255
rect 51 2194 229 2232
rect 269 2221 303 2241
rect 51 2160 85 2194
rect 85 2160 119 2194
rect 119 2160 153 2194
rect 153 2160 187 2194
rect 187 2160 221 2194
rect 221 2160 229 2194
rect 269 2173 296 2182
rect 296 2173 303 2182
rect 51 2122 229 2160
rect 269 2148 303 2173
rect 51 2088 85 2122
rect 85 2088 119 2122
rect 119 2088 153 2122
rect 153 2088 187 2122
rect 187 2088 221 2122
rect 221 2088 229 2122
rect 269 2105 296 2109
rect 296 2105 303 2109
rect 51 2050 229 2088
rect 269 2075 303 2105
rect 51 2016 85 2050
rect 85 2016 119 2050
rect 119 2016 153 2050
rect 153 2016 187 2050
rect 187 2016 221 2050
rect 221 2016 229 2050
rect 51 1978 229 2016
rect 269 2003 303 2036
rect 51 1944 85 1978
rect 85 1944 119 1978
rect 119 1944 153 1978
rect 153 1944 187 1978
rect 187 1944 221 1978
rect 221 1944 229 1978
rect 269 2002 296 2003
rect 296 2002 303 2003
rect 51 1906 229 1944
rect 269 1935 303 1963
rect 51 1872 85 1906
rect 85 1872 119 1906
rect 119 1872 153 1906
rect 153 1872 187 1906
rect 187 1872 221 1906
rect 221 1872 229 1906
rect 269 1929 296 1935
rect 296 1929 303 1935
rect 51 1834 229 1872
rect 269 1867 303 1890
rect 51 1800 85 1834
rect 85 1800 119 1834
rect 119 1800 153 1834
rect 153 1800 187 1834
rect 187 1800 221 1834
rect 221 1800 229 1834
rect 269 1856 296 1867
rect 296 1856 303 1867
rect 51 1762 229 1800
rect 269 1799 303 1817
rect 269 1783 296 1799
rect 296 1783 303 1799
rect 51 1728 85 1762
rect 85 1728 119 1762
rect 119 1728 153 1762
rect 153 1728 187 1762
rect 187 1728 221 1762
rect 221 1728 229 1762
rect 269 1731 303 1744
rect 51 1690 229 1728
rect 269 1710 296 1731
rect 296 1710 303 1731
rect 51 1656 85 1690
rect 85 1656 119 1690
rect 119 1656 153 1690
rect 153 1656 187 1690
rect 187 1656 221 1690
rect 221 1656 229 1690
rect 269 1663 303 1671
rect 51 1618 229 1656
rect 269 1637 296 1663
rect 296 1637 303 1663
rect 51 1584 85 1618
rect 85 1584 119 1618
rect 119 1584 153 1618
rect 153 1584 187 1618
rect 187 1584 221 1618
rect 221 1584 229 1618
rect 269 1595 303 1598
rect 51 1546 229 1584
rect 269 1564 296 1595
rect 296 1564 303 1595
rect 51 1512 85 1546
rect 85 1512 119 1546
rect 119 1512 153 1546
rect 153 1512 187 1546
rect 187 1512 221 1546
rect 221 1512 229 1546
rect 51 1474 229 1512
rect 269 1493 296 1525
rect 296 1493 303 1525
rect 269 1491 303 1493
rect 51 1440 85 1474
rect 85 1440 119 1474
rect 119 1440 153 1474
rect 153 1440 187 1474
rect 187 1440 221 1474
rect 221 1440 229 1474
rect 51 1402 229 1440
rect 269 1425 296 1452
rect 296 1425 303 1452
rect 269 1418 303 1425
rect 51 1368 85 1402
rect 85 1368 119 1402
rect 119 1368 153 1402
rect 153 1368 187 1402
rect 187 1368 221 1402
rect 221 1368 229 1402
rect 51 1330 229 1368
rect 269 1357 296 1379
rect 296 1357 303 1379
rect 269 1345 303 1357
rect 51 1296 85 1330
rect 85 1296 119 1330
rect 119 1296 153 1330
rect 153 1296 187 1330
rect 187 1296 221 1330
rect 221 1296 229 1330
rect 51 1258 229 1296
rect 269 1289 296 1306
rect 296 1289 303 1306
rect 269 1272 303 1289
rect 51 1224 85 1258
rect 85 1224 119 1258
rect 119 1224 153 1258
rect 153 1224 187 1258
rect 187 1224 221 1258
rect 221 1224 229 1258
rect 51 1186 229 1224
rect 269 1221 296 1233
rect 296 1221 303 1233
rect 269 1199 303 1221
rect 51 1152 85 1186
rect 85 1152 119 1186
rect 119 1152 153 1186
rect 153 1152 187 1186
rect 187 1152 221 1186
rect 221 1152 229 1186
rect 269 1153 296 1159
rect 296 1153 303 1159
rect 51 1114 229 1152
rect 269 1125 303 1153
rect 51 1080 85 1114
rect 85 1080 119 1114
rect 119 1080 153 1114
rect 153 1080 187 1114
rect 187 1080 221 1114
rect 221 1080 229 1114
rect 51 1042 229 1080
rect 269 1051 303 1085
rect 51 1008 85 1042
rect 85 1008 119 1042
rect 119 1008 153 1042
rect 153 1008 187 1042
rect 187 1008 221 1042
rect 221 1008 229 1042
rect 51 970 229 1008
rect 269 983 303 1011
rect 51 936 85 970
rect 85 936 119 970
rect 119 936 153 970
rect 153 936 187 970
rect 187 936 221 970
rect 221 936 229 970
rect 269 977 296 983
rect 296 977 303 983
rect 51 898 229 936
rect 269 915 303 937
rect 51 864 85 898
rect 85 864 119 898
rect 119 864 153 898
rect 153 864 187 898
rect 187 864 221 898
rect 221 864 229 898
rect 269 903 296 915
rect 296 903 303 915
rect 51 826 229 864
rect 269 847 303 863
rect 51 792 85 826
rect 85 792 119 826
rect 119 792 153 826
rect 153 792 187 826
rect 187 792 221 826
rect 221 792 229 826
rect 269 829 296 847
rect 296 829 303 847
rect 51 754 229 792
rect 269 779 303 789
rect 51 720 85 754
rect 85 720 119 754
rect 119 720 153 754
rect 153 720 187 754
rect 187 720 221 754
rect 221 720 229 754
rect 269 755 296 779
rect 296 755 303 779
rect 51 682 229 720
rect 269 711 303 715
rect 51 648 85 682
rect 85 648 119 682
rect 119 648 153 682
rect 153 648 187 682
rect 187 648 221 682
rect 221 648 229 682
rect 269 681 296 711
rect 296 681 303 711
rect 51 610 229 648
rect 709 4570 10410 4606
rect 10410 4604 10445 4606
rect 10445 4604 10479 4606
rect 10479 4604 10514 4606
rect 10514 4604 10548 4606
rect 10548 4604 10583 4606
rect 10583 4604 10617 4606
rect 10617 4604 10652 4606
rect 10652 4604 10686 4606
rect 10686 4604 10721 4606
rect 10721 4604 10755 4606
rect 10755 4604 10790 4606
rect 10790 4604 10824 4606
rect 10824 4604 10859 4606
rect 10859 4604 10893 4606
rect 10893 4604 10928 4606
rect 10928 4604 10962 4606
rect 10962 4604 10997 4606
rect 10997 4604 11031 4606
rect 11031 4604 11066 4606
rect 11066 4604 11100 4606
rect 11100 4604 11135 4606
rect 11135 4604 11169 4606
rect 11169 4604 11204 4606
rect 11204 4604 11238 4606
rect 11238 4604 11273 4606
rect 11273 4604 11307 4606
rect 11307 4604 11342 4606
rect 11342 4604 11376 4606
rect 11376 4604 11411 4606
rect 11411 4604 11445 4606
rect 11445 4604 11480 4606
rect 11480 4604 11514 4606
rect 11514 4604 11549 4606
rect 11549 4604 11583 4606
rect 11583 4604 11618 4606
rect 11618 4604 11652 4606
rect 11652 4604 11687 4606
rect 11687 4604 11721 4606
rect 11721 4604 11756 4606
rect 11756 4604 11790 4606
rect 11790 4604 11825 4606
rect 11825 4604 11859 4606
rect 11859 4604 11894 4606
rect 11894 4604 11928 4606
rect 11928 4604 11963 4606
rect 11963 4604 11997 4606
rect 11997 4604 12032 4606
rect 12032 4604 12066 4606
rect 12066 4604 12101 4606
rect 12101 4604 12135 4606
rect 12135 4604 12170 4606
rect 12170 4604 12204 4606
rect 12204 4604 12239 4606
rect 12239 4604 12273 4606
rect 12273 4604 12308 4606
rect 12308 4604 12342 4606
rect 12342 4604 12377 4606
rect 12377 4604 12411 4606
rect 12411 4604 12446 4606
rect 12446 4604 12480 4606
rect 12480 4604 12515 4606
rect 12515 4604 12549 4606
rect 12549 4604 12584 4606
rect 12584 4604 12618 4606
rect 12618 4604 12653 4606
rect 12653 4604 12687 4606
rect 12687 4604 12722 4606
rect 12722 4604 12756 4606
rect 12756 4604 12791 4606
rect 12791 4604 12825 4606
rect 12825 4604 12860 4606
rect 12860 4604 12894 4606
rect 12894 4604 12929 4606
rect 12929 4604 12963 4606
rect 12963 4604 12998 4606
rect 12998 4604 13032 4606
rect 13032 4604 13067 4606
rect 13067 4604 13101 4606
rect 13101 4604 13136 4606
rect 13136 4604 13170 4606
rect 13170 4604 13205 4606
rect 13205 4604 13239 4606
rect 13239 4604 13274 4606
rect 13274 4604 13308 4606
rect 13308 4604 13343 4606
rect 13343 4604 13377 4606
rect 13377 4604 13412 4606
rect 13412 4604 13446 4606
rect 13446 4604 13481 4606
rect 13481 4604 13515 4606
rect 13515 4604 13550 4606
rect 13550 4604 13584 4606
rect 13584 4604 13619 4606
rect 13619 4604 13653 4606
rect 13653 4604 13688 4606
rect 13688 4604 13722 4606
rect 13722 4604 13757 4606
rect 13757 4604 13791 4606
rect 13791 4604 13826 4606
rect 13826 4604 13860 4606
rect 13860 4604 13895 4606
rect 13895 4604 13929 4606
rect 13929 4604 13964 4606
rect 13964 4604 13998 4606
rect 13998 4604 14033 4606
rect 14033 4604 14067 4606
rect 14067 4604 14102 4606
rect 14102 4604 14136 4606
rect 14136 4604 14171 4606
rect 14171 4604 14205 4606
rect 14205 4604 14207 4606
rect 14246 4604 14274 4606
rect 14274 4604 14280 4606
rect 14319 4604 14343 4606
rect 14343 4604 14353 4606
rect 14392 4604 14412 4606
rect 14412 4604 14426 4606
rect 10410 4570 14207 4604
rect 14246 4572 14280 4604
rect 14319 4572 14353 4604
rect 14392 4572 14426 4604
rect 709 4500 12363 4570
rect 12363 4536 12397 4570
rect 12397 4536 12431 4570
rect 12431 4536 12466 4570
rect 12466 4536 12500 4570
rect 12500 4536 12535 4570
rect 12535 4536 12569 4570
rect 12569 4536 12604 4570
rect 12604 4536 12638 4570
rect 12638 4536 12673 4570
rect 12673 4536 12707 4570
rect 12707 4536 12742 4570
rect 12742 4536 12776 4570
rect 12776 4536 12811 4570
rect 12811 4536 12845 4570
rect 12845 4536 12880 4570
rect 12880 4536 12914 4570
rect 12914 4536 12949 4570
rect 12949 4536 12983 4570
rect 12983 4536 13018 4570
rect 13018 4536 13052 4570
rect 13052 4536 13087 4570
rect 13087 4536 13121 4570
rect 13121 4536 13156 4570
rect 13156 4536 13190 4570
rect 13190 4536 13225 4570
rect 13225 4536 13259 4570
rect 13259 4536 13294 4570
rect 13294 4536 13328 4570
rect 13328 4536 13363 4570
rect 13363 4536 13397 4570
rect 13397 4536 13432 4570
rect 13432 4536 13466 4570
rect 13466 4536 13501 4570
rect 13501 4536 13535 4570
rect 13535 4536 13570 4570
rect 13570 4536 13604 4570
rect 13604 4536 13639 4570
rect 13639 4536 13673 4570
rect 13673 4536 13708 4570
rect 13708 4536 13742 4570
rect 13742 4536 13777 4570
rect 13777 4536 13811 4570
rect 13811 4536 13846 4570
rect 13846 4536 13880 4570
rect 13880 4536 13915 4570
rect 13915 4536 13949 4570
rect 13949 4536 13984 4570
rect 13984 4536 14018 4570
rect 14018 4536 14053 4570
rect 14053 4536 14087 4570
rect 14087 4536 14122 4570
rect 14122 4536 14156 4570
rect 14156 4536 14191 4570
rect 14191 4536 14207 4570
rect 12363 4502 14207 4536
rect 14246 4502 14280 4534
rect 14319 4502 14353 4534
rect 14392 4502 14426 4534
rect 12363 4500 12398 4502
rect 12398 4500 12432 4502
rect 12432 4500 12467 4502
rect 12467 4500 12501 4502
rect 12501 4500 12536 4502
rect 12536 4500 12570 4502
rect 12570 4500 12605 4502
rect 12605 4500 12639 4502
rect 12639 4500 12674 4502
rect 12674 4500 12708 4502
rect 12708 4500 12743 4502
rect 12743 4500 12777 4502
rect 12777 4500 12812 4502
rect 12812 4500 12846 4502
rect 12846 4500 12881 4502
rect 12881 4500 12915 4502
rect 12915 4500 12950 4502
rect 12950 4500 12984 4502
rect 12984 4500 13019 4502
rect 13019 4500 13053 4502
rect 13053 4500 13088 4502
rect 13088 4500 13122 4502
rect 13122 4500 13157 4502
rect 13157 4500 13191 4502
rect 13191 4500 13226 4502
rect 13226 4500 13260 4502
rect 13260 4500 13295 4502
rect 13295 4500 13329 4502
rect 13329 4500 13364 4502
rect 13364 4500 13398 4502
rect 13398 4500 13433 4502
rect 13433 4500 13467 4502
rect 13467 4500 13502 4502
rect 13502 4500 13536 4502
rect 13536 4500 13571 4502
rect 13571 4500 13605 4502
rect 13605 4500 13640 4502
rect 13640 4500 13674 4502
rect 13674 4500 13709 4502
rect 13709 4500 13743 4502
rect 13743 4500 13778 4502
rect 13778 4500 13812 4502
rect 13812 4500 13847 4502
rect 13847 4500 13881 4502
rect 13881 4500 13916 4502
rect 13916 4500 13950 4502
rect 13950 4500 13985 4502
rect 13985 4500 14019 4502
rect 14019 4500 14054 4502
rect 14054 4500 14088 4502
rect 14088 4500 14123 4502
rect 14123 4500 14157 4502
rect 14157 4500 14192 4502
rect 14192 4500 14207 4502
rect 14246 4500 14261 4502
rect 14261 4500 14280 4502
rect 14319 4500 14330 4502
rect 14330 4500 14353 4502
rect 14392 4500 14399 4502
rect 14399 4500 14426 4502
rect 674 4445 708 4456
rect 529 4409 563 4426
rect 529 4392 531 4409
rect 531 4392 563 4409
rect 601 4395 633 4426
rect 633 4395 635 4426
rect 601 4392 635 4395
rect 529 4339 563 4351
rect 529 4317 531 4339
rect 531 4317 563 4339
rect 601 4322 633 4351
rect 633 4322 635 4351
rect 601 4317 635 4322
rect 529 4269 563 4276
rect 529 4242 531 4269
rect 531 4242 563 4269
rect 601 4249 633 4276
rect 633 4249 635 4276
rect 601 4242 635 4249
rect 529 4199 563 4201
rect 529 4167 531 4199
rect 531 4167 563 4199
rect 601 4177 633 4201
rect 633 4177 635 4201
rect 601 4167 635 4177
rect 529 4095 531 4126
rect 531 4095 563 4126
rect 601 4105 633 4126
rect 633 4105 635 4126
rect 529 4092 563 4095
rect 601 4092 635 4105
rect 674 4082 780 4445
rect 14356 4398 14390 4432
rect 14428 4426 14462 4456
rect 14356 4325 14390 4359
rect 529 4025 531 4052
rect 531 4025 563 4052
rect 601 4033 633 4052
rect 633 4033 635 4052
rect 674 4048 745 4082
rect 745 4048 779 4082
rect 779 4048 780 4082
rect 529 4018 563 4025
rect 601 4018 635 4033
rect 674 4014 780 4048
rect 529 3955 531 3978
rect 531 3955 563 3978
rect 601 3961 633 3978
rect 633 3961 635 3978
rect 674 3980 745 4014
rect 745 3980 779 4014
rect 779 3980 780 4014
rect 529 3944 563 3955
rect 601 3944 635 3961
rect 674 3946 780 3980
rect 529 3886 531 3904
rect 531 3886 563 3904
rect 601 3889 633 3904
rect 633 3889 635 3904
rect 674 3912 745 3946
rect 745 3912 779 3946
rect 779 3912 780 3946
rect 529 3870 563 3886
rect 601 3870 635 3889
rect 674 3878 780 3912
rect 674 3844 745 3878
rect 745 3844 779 3878
rect 779 3844 780 3878
rect 674 3810 780 3844
rect 529 3760 563 3794
rect 601 3760 635 3794
rect 674 3776 745 3810
rect 745 3776 779 3810
rect 779 3776 780 3810
rect 529 3715 531 3720
rect 531 3715 563 3720
rect 601 3715 633 3720
rect 633 3715 635 3720
rect 674 3742 780 3776
rect 529 3686 563 3715
rect 601 3686 635 3715
rect 674 3708 745 3742
rect 745 3708 779 3742
rect 779 3708 780 3742
rect 674 3674 780 3708
rect 529 3612 563 3646
rect 601 3612 635 3646
rect 674 3640 745 3674
rect 745 3640 779 3674
rect 779 3640 780 3674
rect 674 3606 780 3640
rect 674 3572 745 3606
rect 745 3572 779 3606
rect 779 3572 780 3606
rect 529 3542 563 3572
rect 601 3542 635 3572
rect 529 3538 531 3542
rect 531 3538 563 3542
rect 601 3538 633 3542
rect 633 3538 635 3542
rect 674 3538 780 3572
rect 674 3504 745 3538
rect 745 3504 779 3538
rect 779 3504 780 3538
rect 529 3473 563 3498
rect 601 3473 635 3498
rect 529 3464 531 3473
rect 531 3464 563 3473
rect 601 3464 633 3473
rect 633 3464 635 3473
rect 674 3470 780 3504
rect 674 3436 745 3470
rect 745 3436 779 3470
rect 779 3436 780 3470
rect 529 3404 563 3424
rect 601 3404 635 3424
rect 529 3390 531 3404
rect 531 3390 563 3404
rect 601 3390 633 3404
rect 633 3390 635 3404
rect 674 3402 780 3436
rect 674 3368 745 3402
rect 745 3368 779 3402
rect 779 3368 780 3402
rect 529 3335 563 3350
rect 601 3335 635 3350
rect 529 3316 531 3335
rect 531 3316 563 3335
rect 601 3316 633 3335
rect 633 3316 635 3335
rect 674 3334 780 3368
rect 674 3300 745 3334
rect 745 3300 779 3334
rect 779 3300 780 3334
rect 529 3266 563 3276
rect 601 3266 635 3276
rect 674 3266 780 3300
rect 529 3242 531 3266
rect 531 3242 563 3266
rect 601 3242 633 3266
rect 633 3242 635 3266
rect 674 3232 745 3266
rect 745 3232 779 3266
rect 779 3232 780 3266
rect 529 3197 563 3202
rect 601 3197 635 3202
rect 674 3198 780 3232
rect 529 3168 531 3197
rect 531 3168 563 3197
rect 601 3168 633 3197
rect 633 3168 635 3197
rect 674 3164 745 3198
rect 745 3164 779 3198
rect 779 3164 780 3198
rect 529 3094 531 3128
rect 531 3094 563 3128
rect 601 3094 633 3128
rect 633 3094 635 3128
rect 529 3025 531 3054
rect 531 3025 563 3054
rect 601 3025 633 3054
rect 633 3025 635 3054
rect 529 3020 563 3025
rect 601 3020 635 3025
rect 529 2956 531 2980
rect 531 2956 563 2980
rect 601 2956 633 2980
rect 633 2956 635 2980
rect 529 2946 563 2956
rect 601 2946 635 2956
rect 529 2887 531 2906
rect 531 2887 563 2906
rect 601 2887 633 2906
rect 633 2887 635 2906
rect 529 2872 563 2887
rect 601 2872 635 2887
rect 529 2818 531 2832
rect 531 2818 563 2832
rect 601 2818 633 2832
rect 633 2818 635 2832
rect 529 2798 563 2818
rect 601 2798 635 2818
rect 529 2749 531 2758
rect 531 2749 563 2758
rect 601 2749 633 2758
rect 633 2749 635 2758
rect 529 2724 563 2749
rect 601 2724 635 2749
rect 529 2680 531 2684
rect 531 2680 563 2684
rect 601 2680 633 2684
rect 633 2680 635 2684
rect 529 2650 563 2680
rect 601 2650 635 2680
rect 529 2576 563 2610
rect 601 2576 635 2610
rect 529 2507 563 2536
rect 601 2507 635 2536
rect 529 2502 531 2507
rect 531 2502 563 2507
rect 601 2502 633 2507
rect 633 2502 635 2507
rect 674 2482 780 3164
rect 529 2438 563 2462
rect 601 2438 635 2462
rect 674 2448 745 2482
rect 745 2448 779 2482
rect 779 2448 780 2482
rect 529 2428 531 2438
rect 531 2428 563 2438
rect 601 2428 633 2438
rect 633 2428 635 2438
rect 674 2414 780 2448
rect 529 2369 563 2389
rect 601 2369 635 2389
rect 674 2380 745 2414
rect 745 2380 779 2414
rect 779 2380 780 2414
rect 529 2355 531 2369
rect 531 2355 563 2369
rect 601 2355 633 2369
rect 633 2355 635 2369
rect 674 2346 780 2380
rect 529 2300 563 2316
rect 601 2300 635 2316
rect 674 2312 745 2346
rect 745 2312 779 2346
rect 779 2312 780 2346
rect 529 2282 531 2300
rect 531 2282 563 2300
rect 601 2282 633 2300
rect 633 2282 635 2300
rect 674 2278 780 2312
rect 674 2244 745 2278
rect 745 2244 779 2278
rect 779 2244 780 2278
rect 529 2231 563 2243
rect 601 2231 635 2243
rect 529 2209 531 2231
rect 531 2209 563 2231
rect 601 2209 633 2231
rect 633 2209 635 2231
rect 674 2210 780 2244
rect 674 2176 745 2210
rect 745 2176 779 2210
rect 779 2176 780 2210
rect 529 2163 563 2170
rect 529 2136 531 2163
rect 531 2136 563 2163
rect 601 2162 635 2170
rect 601 2136 633 2162
rect 633 2136 635 2162
rect 674 2142 780 2176
rect 674 2108 745 2142
rect 745 2108 779 2142
rect 779 2108 780 2142
rect 529 2095 563 2097
rect 529 2063 531 2095
rect 531 2063 563 2095
rect 601 2093 635 2097
rect 601 2063 633 2093
rect 633 2063 635 2093
rect 674 2074 780 2108
rect 674 2040 745 2074
rect 745 2040 779 2074
rect 779 2040 780 2074
rect 529 1993 531 2024
rect 531 1993 563 2024
rect 529 1990 563 1993
rect 601 1990 633 2024
rect 633 1990 635 2024
rect 674 2006 780 2040
rect 674 1972 745 2006
rect 745 1972 779 2006
rect 779 1972 780 2006
rect 529 1925 531 1951
rect 531 1925 563 1951
rect 529 1917 563 1925
rect 601 1921 633 1951
rect 633 1921 635 1951
rect 674 1938 780 1972
rect 601 1917 635 1921
rect 674 1904 745 1938
rect 745 1904 779 1938
rect 779 1904 780 1938
rect 529 1857 531 1878
rect 531 1857 563 1878
rect 529 1844 563 1857
rect 601 1852 633 1878
rect 633 1852 635 1878
rect 674 1870 780 1904
rect 601 1844 635 1852
rect 674 1836 745 1870
rect 745 1836 779 1870
rect 779 1836 780 1870
rect 529 1789 531 1805
rect 531 1789 563 1805
rect 529 1771 563 1789
rect 601 1783 633 1805
rect 633 1783 635 1805
rect 674 1802 780 1836
rect 601 1771 635 1783
rect 674 1768 745 1802
rect 745 1768 779 1802
rect 779 1768 780 1802
rect 529 1721 531 1732
rect 531 1721 563 1732
rect 529 1698 563 1721
rect 601 1714 633 1732
rect 633 1714 635 1732
rect 674 1734 780 1768
rect 601 1698 635 1714
rect 674 1700 745 1734
rect 745 1700 779 1734
rect 779 1700 780 1734
rect 529 1653 531 1659
rect 531 1653 563 1659
rect 529 1625 563 1653
rect 601 1645 633 1659
rect 633 1645 635 1659
rect 674 1666 780 1700
rect 601 1625 635 1645
rect 674 1632 745 1666
rect 745 1632 779 1666
rect 779 1632 780 1666
rect 529 1585 531 1586
rect 531 1585 563 1586
rect 529 1552 563 1585
rect 601 1576 633 1586
rect 633 1576 635 1586
rect 674 1598 780 1632
rect 601 1552 635 1576
rect 674 1564 745 1598
rect 745 1564 779 1598
rect 779 1564 780 1598
rect 529 1483 563 1513
rect 601 1507 633 1513
rect 633 1507 635 1513
rect 529 1479 531 1483
rect 531 1479 563 1483
rect 601 1479 635 1507
rect 529 1415 563 1440
rect 601 1438 633 1440
rect 633 1438 635 1440
rect 529 1406 531 1415
rect 531 1406 563 1415
rect 601 1406 635 1438
rect 529 1347 563 1367
rect 529 1333 531 1347
rect 531 1333 563 1347
rect 601 1334 635 1367
rect 601 1333 633 1334
rect 633 1333 635 1334
rect 529 1279 563 1294
rect 529 1260 531 1279
rect 531 1260 563 1279
rect 601 1265 635 1294
rect 601 1260 633 1265
rect 633 1260 635 1265
rect 529 1211 563 1221
rect 529 1187 531 1211
rect 531 1187 563 1211
rect 601 1196 635 1221
rect 601 1187 633 1196
rect 633 1187 635 1196
rect 529 1143 563 1148
rect 529 1114 531 1143
rect 531 1114 563 1143
rect 601 1127 635 1148
rect 601 1114 633 1127
rect 633 1114 635 1127
rect 529 1041 531 1075
rect 531 1041 563 1075
rect 601 1058 635 1075
rect 601 1041 633 1058
rect 633 1041 635 1058
rect 529 973 531 1002
rect 531 973 563 1002
rect 601 989 635 1002
rect 529 968 563 973
rect 601 968 633 989
rect 633 968 635 989
rect 529 920 531 929
rect 531 920 563 929
rect 601 920 635 929
rect 529 895 563 920
rect 601 895 635 920
rect 674 894 780 1564
rect 1067 4064 1101 4098
rect 1139 4064 1173 4098
rect 1211 4064 1245 4098
rect 1067 3991 1101 4025
rect 1139 3991 1173 4025
rect 1211 3991 1245 4025
rect 1067 3918 1101 3952
rect 1139 3918 1173 3952
rect 1211 3918 1245 3952
rect 1067 3845 1101 3879
rect 1139 3845 1173 3879
rect 1211 3845 1245 3879
rect 1067 3772 1101 3806
rect 1139 3772 1173 3806
rect 1211 3772 1245 3806
rect 1067 3699 1101 3733
rect 1139 3699 1173 3733
rect 1211 3699 1245 3733
rect 1067 3626 1101 3660
rect 1139 3626 1173 3660
rect 1211 3626 1245 3660
rect 1067 3553 1101 3587
rect 1139 3553 1173 3587
rect 1211 3553 1245 3587
rect 1067 3480 1101 3514
rect 1139 3480 1173 3514
rect 1211 3480 1245 3514
rect 1067 3407 1101 3441
rect 1139 3407 1173 3441
rect 1211 3407 1245 3441
rect 1067 3334 1101 3368
rect 1139 3334 1173 3368
rect 1211 3334 1245 3368
rect 1067 3261 1101 3295
rect 1139 3261 1173 3295
rect 1211 3261 1245 3295
rect 1067 3188 1101 3222
rect 1139 3188 1173 3222
rect 1211 3188 1245 3222
rect 1067 3115 1101 3149
rect 1139 3115 1173 3149
rect 1211 3115 1245 3149
rect 1067 3042 1101 3076
rect 1139 3042 1173 3076
rect 1211 3042 1245 3076
rect 1067 2969 1101 3003
rect 1139 2969 1173 3003
rect 1211 2969 1245 3003
rect 1067 2896 1101 2930
rect 1139 2896 1173 2930
rect 1211 2896 1245 2930
rect 1067 2823 1101 2857
rect 1139 2823 1173 2857
rect 1211 2823 1245 2857
rect 1067 2750 1101 2784
rect 1139 2750 1173 2784
rect 1211 2750 1245 2784
rect 1067 2677 1101 2711
rect 1139 2677 1173 2711
rect 1211 2677 1245 2711
rect 1067 2604 1101 2638
rect 1139 2604 1173 2638
rect 1211 2604 1245 2638
rect 1067 2531 1101 2565
rect 1139 2531 1173 2565
rect 1211 2531 1245 2565
rect 1067 2458 1101 2492
rect 1139 2458 1173 2492
rect 1211 2458 1245 2492
rect 1067 2385 1101 2419
rect 1139 2385 1173 2419
rect 1211 2385 1245 2419
rect 1067 2312 1101 2346
rect 1139 2312 1173 2346
rect 1211 2312 1245 2346
rect 1067 2239 1101 2273
rect 1139 2239 1173 2273
rect 1211 2239 1245 2273
rect 1067 2166 1101 2200
rect 1139 2166 1173 2200
rect 1211 2166 1245 2200
rect 1067 2092 1101 2126
rect 1139 2092 1173 2126
rect 1211 2092 1245 2126
rect 1067 2018 1101 2052
rect 1139 2018 1173 2052
rect 1211 2018 1245 2052
rect 1067 1944 1101 1978
rect 1139 1944 1173 1978
rect 1211 1944 1245 1978
rect 1067 1870 1101 1904
rect 1139 1870 1173 1904
rect 1211 1870 1245 1904
rect 1067 1796 1101 1830
rect 1139 1796 1173 1830
rect 1211 1796 1245 1830
rect 1067 1722 1101 1756
rect 1139 1722 1173 1756
rect 1211 1722 1245 1756
rect 1067 1648 1101 1682
rect 1139 1648 1173 1682
rect 1211 1648 1245 1682
rect 1067 1574 1101 1608
rect 1139 1574 1173 1608
rect 1211 1574 1245 1608
rect 924 1216 958 1250
rect 924 1144 958 1178
rect 1635 4092 1669 4118
rect 1563 4082 1741 4092
rect 1563 4048 1567 4082
rect 1567 4048 1635 4082
rect 1635 4048 1669 4082
rect 1669 4048 1737 4082
rect 1737 4048 1741 4082
rect 1563 4014 1741 4048
rect 1563 3980 1567 4014
rect 1567 3980 1635 4014
rect 1635 3980 1669 4014
rect 1669 3980 1737 4014
rect 1737 3980 1741 4014
rect 1563 3946 1741 3980
rect 1563 3912 1567 3946
rect 1567 3912 1635 3946
rect 1635 3912 1669 3946
rect 1669 3912 1737 3946
rect 1737 3912 1741 3946
rect 1563 3878 1741 3912
rect 1563 3844 1567 3878
rect 1567 3844 1635 3878
rect 1635 3844 1669 3878
rect 1669 3844 1737 3878
rect 1737 3844 1741 3878
rect 1563 3810 1741 3844
rect 1563 3776 1567 3810
rect 1567 3776 1635 3810
rect 1635 3776 1669 3810
rect 1669 3776 1737 3810
rect 1737 3776 1741 3810
rect 1563 3742 1741 3776
rect 1563 3708 1567 3742
rect 1567 3708 1635 3742
rect 1635 3708 1669 3742
rect 1669 3708 1737 3742
rect 1737 3708 1741 3742
rect 1563 3674 1741 3708
rect 1563 3640 1567 3674
rect 1567 3640 1635 3674
rect 1635 3640 1669 3674
rect 1669 3640 1737 3674
rect 1737 3640 1741 3674
rect 1563 3606 1741 3640
rect 1563 3572 1567 3606
rect 1567 3572 1635 3606
rect 1635 3572 1669 3606
rect 1669 3572 1737 3606
rect 1737 3572 1741 3606
rect 1563 3538 1741 3572
rect 1563 3504 1567 3538
rect 1567 3504 1635 3538
rect 1635 3504 1669 3538
rect 1669 3504 1737 3538
rect 1737 3504 1741 3538
rect 1563 3470 1741 3504
rect 1563 3436 1567 3470
rect 1567 3436 1635 3470
rect 1635 3436 1669 3470
rect 1669 3436 1737 3470
rect 1737 3436 1741 3470
rect 1563 3402 1741 3436
rect 1563 3368 1567 3402
rect 1567 3368 1635 3402
rect 1635 3368 1669 3402
rect 1669 3368 1737 3402
rect 1737 3368 1741 3402
rect 1563 3334 1741 3368
rect 1563 3300 1567 3334
rect 1567 3300 1635 3334
rect 1635 3300 1669 3334
rect 1669 3300 1737 3334
rect 1737 3300 1741 3334
rect 1563 3266 1741 3300
rect 1563 3232 1567 3266
rect 1567 3232 1635 3266
rect 1635 3232 1669 3266
rect 1669 3232 1737 3266
rect 1737 3232 1741 3266
rect 1563 3198 1741 3232
rect 1563 3194 1567 3198
rect 1567 3194 1635 3198
rect 1635 3194 1669 3198
rect 1669 3194 1737 3198
rect 1737 3194 1741 3198
rect 1635 3164 1669 3182
rect 1635 3148 1669 3164
rect 1563 3074 1597 3108
rect 1635 3074 1669 3108
rect 1707 3074 1741 3108
rect 1563 2994 1597 3028
rect 1635 2994 1669 3028
rect 1707 2994 1741 3028
rect 1563 2914 1597 2948
rect 1635 2914 1669 2948
rect 1707 2914 1741 2948
rect 1563 2834 1597 2868
rect 1635 2834 1669 2868
rect 1707 2834 1741 2868
rect 1563 2754 1597 2788
rect 1635 2754 1669 2788
rect 1707 2754 1741 2788
rect 1563 2674 1597 2708
rect 1635 2674 1669 2708
rect 1707 2674 1741 2708
rect 1563 2594 1597 2628
rect 1635 2594 1669 2628
rect 1707 2594 1741 2628
rect 1635 2540 1669 2556
rect 1635 2522 1669 2540
rect 1563 2506 1567 2518
rect 1567 2506 1635 2518
rect 1635 2506 1669 2518
rect 1669 2506 1737 2518
rect 1737 2506 1741 2518
rect 1563 2472 1741 2506
rect 1563 2438 1567 2472
rect 1567 2438 1635 2472
rect 1635 2438 1669 2472
rect 1669 2438 1737 2472
rect 1737 2438 1741 2472
rect 1563 2404 1741 2438
rect 1563 2370 1567 2404
rect 1567 2370 1635 2404
rect 1635 2370 1669 2404
rect 1669 2370 1737 2404
rect 1737 2370 1741 2404
rect 1563 2336 1741 2370
rect 1563 2302 1567 2336
rect 1567 2302 1635 2336
rect 1635 2302 1669 2336
rect 1669 2302 1737 2336
rect 1737 2302 1741 2336
rect 1563 2268 1741 2302
rect 1563 2234 1567 2268
rect 1567 2234 1635 2268
rect 1635 2234 1669 2268
rect 1669 2234 1737 2268
rect 1737 2234 1741 2268
rect 1563 2200 1741 2234
rect 1563 2166 1567 2200
rect 1567 2166 1635 2200
rect 1635 2166 1669 2200
rect 1669 2166 1737 2200
rect 1737 2166 1741 2200
rect 1563 2132 1741 2166
rect 1563 2098 1567 2132
rect 1567 2098 1635 2132
rect 1635 2098 1669 2132
rect 1669 2098 1737 2132
rect 1737 2098 1741 2132
rect 1563 2064 1741 2098
rect 1563 2030 1567 2064
rect 1567 2030 1635 2064
rect 1635 2030 1669 2064
rect 1669 2030 1737 2064
rect 1737 2030 1741 2064
rect 1563 1996 1741 2030
rect 1563 1962 1567 1996
rect 1567 1962 1635 1996
rect 1635 1962 1669 1996
rect 1669 1962 1737 1996
rect 1737 1962 1741 1996
rect 1563 1928 1741 1962
rect 1563 1894 1567 1928
rect 1567 1894 1635 1928
rect 1635 1894 1669 1928
rect 1669 1894 1737 1928
rect 1737 1894 1741 1928
rect 1563 1860 1741 1894
rect 1563 1826 1567 1860
rect 1567 1826 1635 1860
rect 1635 1826 1669 1860
rect 1669 1826 1737 1860
rect 1737 1826 1741 1860
rect 1563 1792 1741 1826
rect 1563 1758 1567 1792
rect 1567 1758 1635 1792
rect 1635 1758 1669 1792
rect 1669 1758 1737 1792
rect 1737 1758 1741 1792
rect 1563 1724 1741 1758
rect 1563 1690 1567 1724
rect 1567 1690 1635 1724
rect 1635 1690 1669 1724
rect 1669 1690 1737 1724
rect 1737 1690 1741 1724
rect 1563 1656 1741 1690
rect 1563 1622 1567 1656
rect 1567 1622 1635 1656
rect 1635 1622 1669 1656
rect 1669 1622 1737 1656
rect 1737 1622 1741 1656
rect 1563 1620 1741 1622
rect 1635 1586 1669 1620
rect 1318 1144 1424 1250
rect 2059 4064 2093 4098
rect 2131 4064 2165 4098
rect 2203 4064 2237 4098
rect 2059 3991 2093 4025
rect 2131 3991 2165 4025
rect 2203 3991 2237 4025
rect 2059 3918 2093 3952
rect 2131 3918 2165 3952
rect 2203 3918 2237 3952
rect 2059 3845 2093 3879
rect 2131 3845 2165 3879
rect 2203 3845 2237 3879
rect 2059 3772 2093 3806
rect 2131 3772 2165 3806
rect 2203 3772 2237 3806
rect 2059 3699 2093 3733
rect 2131 3699 2165 3733
rect 2203 3699 2237 3733
rect 2059 3626 2093 3660
rect 2131 3626 2165 3660
rect 2203 3626 2237 3660
rect 2059 3553 2093 3587
rect 2131 3553 2165 3587
rect 2203 3553 2237 3587
rect 2059 3480 2093 3514
rect 2131 3480 2165 3514
rect 2203 3480 2237 3514
rect 2059 3407 2093 3441
rect 2131 3407 2165 3441
rect 2203 3407 2237 3441
rect 2059 3334 2093 3368
rect 2131 3334 2165 3368
rect 2203 3334 2237 3368
rect 2059 3261 2093 3295
rect 2131 3261 2165 3295
rect 2203 3261 2237 3295
rect 2059 3188 2093 3222
rect 2131 3188 2165 3222
rect 2203 3188 2237 3222
rect 2059 3115 2093 3149
rect 2131 3115 2165 3149
rect 2203 3115 2237 3149
rect 2059 3042 2093 3076
rect 2131 3042 2165 3076
rect 2203 3042 2237 3076
rect 2059 2969 2093 3003
rect 2131 2969 2165 3003
rect 2203 2969 2237 3003
rect 2059 2896 2093 2930
rect 2131 2896 2165 2930
rect 2203 2896 2237 2930
rect 2059 2823 2093 2857
rect 2131 2823 2165 2857
rect 2203 2823 2237 2857
rect 2059 2750 2093 2784
rect 2131 2750 2165 2784
rect 2203 2750 2237 2784
rect 2059 2677 2093 2711
rect 2131 2677 2165 2711
rect 2203 2677 2237 2711
rect 2059 2604 2093 2638
rect 2131 2604 2165 2638
rect 2203 2604 2237 2638
rect 2059 2531 2093 2565
rect 2131 2531 2165 2565
rect 2203 2531 2237 2565
rect 2059 2458 2093 2492
rect 2131 2458 2165 2492
rect 2203 2458 2237 2492
rect 2059 2385 2093 2419
rect 2131 2385 2165 2419
rect 2203 2385 2237 2419
rect 2059 2312 2093 2346
rect 2131 2312 2165 2346
rect 2203 2312 2237 2346
rect 2059 2239 2093 2273
rect 2131 2239 2165 2273
rect 2203 2239 2237 2273
rect 2059 2166 2093 2200
rect 2131 2166 2165 2200
rect 2203 2166 2237 2200
rect 2059 2092 2093 2126
rect 2131 2092 2165 2126
rect 2203 2092 2237 2126
rect 2059 2018 2093 2052
rect 2131 2018 2165 2052
rect 2203 2018 2237 2052
rect 2059 1944 2093 1978
rect 2131 1944 2165 1978
rect 2203 1944 2237 1978
rect 2059 1870 2093 1904
rect 2131 1870 2165 1904
rect 2203 1870 2237 1904
rect 2059 1796 2093 1830
rect 2131 1796 2165 1830
rect 2203 1796 2237 1830
rect 2059 1722 2093 1756
rect 2131 1722 2165 1756
rect 2203 1722 2237 1756
rect 2059 1648 2093 1682
rect 2131 1648 2165 1682
rect 2203 1648 2237 1682
rect 2059 1574 2093 1608
rect 2131 1574 2165 1608
rect 2203 1574 2237 1608
rect 1880 1144 1986 1250
rect 2627 4092 2661 4118
rect 2555 4082 2733 4092
rect 2555 4048 2559 4082
rect 2559 4048 2627 4082
rect 2627 4048 2661 4082
rect 2661 4048 2729 4082
rect 2729 4048 2733 4082
rect 2555 4014 2733 4048
rect 2555 3980 2559 4014
rect 2559 3980 2627 4014
rect 2627 3980 2661 4014
rect 2661 3980 2729 4014
rect 2729 3980 2733 4014
rect 2555 3946 2733 3980
rect 2555 3912 2559 3946
rect 2559 3912 2627 3946
rect 2627 3912 2661 3946
rect 2661 3912 2729 3946
rect 2729 3912 2733 3946
rect 2555 3878 2733 3912
rect 2555 3844 2559 3878
rect 2559 3844 2627 3878
rect 2627 3844 2661 3878
rect 2661 3844 2729 3878
rect 2729 3844 2733 3878
rect 2555 3810 2733 3844
rect 2555 3776 2559 3810
rect 2559 3776 2627 3810
rect 2627 3776 2661 3810
rect 2661 3776 2729 3810
rect 2729 3776 2733 3810
rect 2555 3742 2733 3776
rect 2555 3708 2559 3742
rect 2559 3708 2627 3742
rect 2627 3708 2661 3742
rect 2661 3708 2729 3742
rect 2729 3708 2733 3742
rect 2555 3674 2733 3708
rect 2555 3640 2559 3674
rect 2559 3640 2627 3674
rect 2627 3640 2661 3674
rect 2661 3640 2729 3674
rect 2729 3640 2733 3674
rect 2555 3606 2733 3640
rect 2555 3572 2559 3606
rect 2559 3572 2627 3606
rect 2627 3572 2661 3606
rect 2661 3572 2729 3606
rect 2729 3572 2733 3606
rect 2555 3538 2733 3572
rect 2555 3504 2559 3538
rect 2559 3504 2627 3538
rect 2627 3504 2661 3538
rect 2661 3504 2729 3538
rect 2729 3504 2733 3538
rect 2555 3470 2733 3504
rect 2555 3436 2559 3470
rect 2559 3436 2627 3470
rect 2627 3436 2661 3470
rect 2661 3436 2729 3470
rect 2729 3436 2733 3470
rect 2555 3402 2733 3436
rect 2555 3368 2559 3402
rect 2559 3368 2627 3402
rect 2627 3368 2661 3402
rect 2661 3368 2729 3402
rect 2729 3368 2733 3402
rect 2555 3334 2733 3368
rect 2555 3300 2559 3334
rect 2559 3300 2627 3334
rect 2627 3300 2661 3334
rect 2661 3300 2729 3334
rect 2729 3300 2733 3334
rect 2555 3266 2733 3300
rect 2555 3232 2559 3266
rect 2559 3232 2627 3266
rect 2627 3232 2661 3266
rect 2661 3232 2729 3266
rect 2729 3232 2733 3266
rect 2555 3198 2733 3232
rect 2555 3194 2559 3198
rect 2559 3194 2627 3198
rect 2627 3194 2661 3198
rect 2661 3194 2729 3198
rect 2729 3194 2733 3198
rect 2627 3164 2661 3182
rect 2627 3148 2661 3164
rect 2555 3074 2589 3108
rect 2627 3074 2661 3108
rect 2699 3074 2733 3108
rect 2555 2994 2589 3028
rect 2627 2994 2661 3028
rect 2699 2994 2733 3028
rect 2555 2914 2589 2948
rect 2627 2914 2661 2948
rect 2699 2914 2733 2948
rect 2555 2834 2589 2868
rect 2627 2834 2661 2868
rect 2699 2834 2733 2868
rect 2555 2754 2589 2788
rect 2627 2754 2661 2788
rect 2699 2754 2733 2788
rect 2555 2674 2589 2708
rect 2627 2674 2661 2708
rect 2699 2674 2733 2708
rect 2555 2594 2589 2628
rect 2627 2594 2661 2628
rect 2699 2594 2733 2628
rect 2627 2540 2661 2556
rect 2627 2522 2661 2540
rect 2555 2506 2559 2518
rect 2559 2506 2627 2518
rect 2627 2506 2661 2518
rect 2661 2506 2729 2518
rect 2729 2506 2733 2518
rect 2555 2472 2733 2506
rect 2555 2438 2559 2472
rect 2559 2438 2627 2472
rect 2627 2438 2661 2472
rect 2661 2438 2729 2472
rect 2729 2438 2733 2472
rect 2555 2404 2733 2438
rect 2555 2370 2559 2404
rect 2559 2370 2627 2404
rect 2627 2370 2661 2404
rect 2661 2370 2729 2404
rect 2729 2370 2733 2404
rect 2555 2336 2733 2370
rect 2555 2302 2559 2336
rect 2559 2302 2627 2336
rect 2627 2302 2661 2336
rect 2661 2302 2729 2336
rect 2729 2302 2733 2336
rect 2555 2268 2733 2302
rect 2555 2234 2559 2268
rect 2559 2234 2627 2268
rect 2627 2234 2661 2268
rect 2661 2234 2729 2268
rect 2729 2234 2733 2268
rect 2555 2200 2733 2234
rect 2555 2166 2559 2200
rect 2559 2166 2627 2200
rect 2627 2166 2661 2200
rect 2661 2166 2729 2200
rect 2729 2166 2733 2200
rect 2555 2132 2733 2166
rect 2555 2098 2559 2132
rect 2559 2098 2627 2132
rect 2627 2098 2661 2132
rect 2661 2098 2729 2132
rect 2729 2098 2733 2132
rect 2555 2064 2733 2098
rect 2555 2030 2559 2064
rect 2559 2030 2627 2064
rect 2627 2030 2661 2064
rect 2661 2030 2729 2064
rect 2729 2030 2733 2064
rect 2555 1996 2733 2030
rect 2555 1962 2559 1996
rect 2559 1962 2627 1996
rect 2627 1962 2661 1996
rect 2661 1962 2729 1996
rect 2729 1962 2733 1996
rect 2555 1928 2733 1962
rect 2555 1894 2559 1928
rect 2559 1894 2627 1928
rect 2627 1894 2661 1928
rect 2661 1894 2729 1928
rect 2729 1894 2733 1928
rect 2555 1860 2733 1894
rect 2555 1826 2559 1860
rect 2559 1826 2627 1860
rect 2627 1826 2661 1860
rect 2661 1826 2729 1860
rect 2729 1826 2733 1860
rect 2555 1792 2733 1826
rect 2555 1758 2559 1792
rect 2559 1758 2627 1792
rect 2627 1758 2661 1792
rect 2661 1758 2729 1792
rect 2729 1758 2733 1792
rect 2555 1724 2733 1758
rect 2555 1690 2559 1724
rect 2559 1690 2627 1724
rect 2627 1690 2661 1724
rect 2661 1690 2729 1724
rect 2729 1690 2733 1724
rect 2555 1656 2733 1690
rect 2555 1622 2559 1656
rect 2559 1622 2627 1656
rect 2627 1622 2661 1656
rect 2661 1622 2729 1656
rect 2729 1622 2733 1656
rect 2555 1620 2733 1622
rect 2627 1586 2661 1620
rect 2310 1144 2416 1250
rect 3051 4064 3085 4098
rect 3123 4064 3157 4098
rect 3195 4064 3229 4098
rect 3051 3991 3085 4025
rect 3123 3991 3157 4025
rect 3195 3991 3229 4025
rect 3051 3918 3085 3952
rect 3123 3918 3157 3952
rect 3195 3918 3229 3952
rect 3051 3845 3085 3879
rect 3123 3845 3157 3879
rect 3195 3845 3229 3879
rect 3051 3772 3085 3806
rect 3123 3772 3157 3806
rect 3195 3772 3229 3806
rect 3051 3699 3085 3733
rect 3123 3699 3157 3733
rect 3195 3699 3229 3733
rect 3051 3626 3085 3660
rect 3123 3626 3157 3660
rect 3195 3626 3229 3660
rect 3051 3553 3085 3587
rect 3123 3553 3157 3587
rect 3195 3553 3229 3587
rect 3051 3480 3085 3514
rect 3123 3480 3157 3514
rect 3195 3480 3229 3514
rect 3051 3407 3085 3441
rect 3123 3407 3157 3441
rect 3195 3407 3229 3441
rect 3051 3334 3085 3368
rect 3123 3334 3157 3368
rect 3195 3334 3229 3368
rect 3051 3261 3085 3295
rect 3123 3261 3157 3295
rect 3195 3261 3229 3295
rect 3051 3188 3085 3222
rect 3123 3188 3157 3222
rect 3195 3188 3229 3222
rect 3051 3115 3085 3149
rect 3123 3115 3157 3149
rect 3195 3115 3229 3149
rect 3051 3042 3085 3076
rect 3123 3042 3157 3076
rect 3195 3042 3229 3076
rect 3051 2969 3085 3003
rect 3123 2969 3157 3003
rect 3195 2969 3229 3003
rect 3051 2896 3085 2930
rect 3123 2896 3157 2930
rect 3195 2896 3229 2930
rect 3051 2823 3085 2857
rect 3123 2823 3157 2857
rect 3195 2823 3229 2857
rect 3051 2750 3085 2784
rect 3123 2750 3157 2784
rect 3195 2750 3229 2784
rect 3051 2677 3085 2711
rect 3123 2677 3157 2711
rect 3195 2677 3229 2711
rect 3051 2604 3085 2638
rect 3123 2604 3157 2638
rect 3195 2604 3229 2638
rect 3051 2531 3085 2565
rect 3123 2531 3157 2565
rect 3195 2531 3229 2565
rect 3051 2458 3085 2492
rect 3123 2458 3157 2492
rect 3195 2458 3229 2492
rect 3051 2385 3085 2419
rect 3123 2385 3157 2419
rect 3195 2385 3229 2419
rect 3051 2312 3085 2346
rect 3123 2312 3157 2346
rect 3195 2312 3229 2346
rect 3051 2239 3085 2273
rect 3123 2239 3157 2273
rect 3195 2239 3229 2273
rect 3051 2166 3085 2200
rect 3123 2166 3157 2200
rect 3195 2166 3229 2200
rect 3051 2092 3085 2126
rect 3123 2092 3157 2126
rect 3195 2092 3229 2126
rect 3051 2018 3085 2052
rect 3123 2018 3157 2052
rect 3195 2018 3229 2052
rect 3051 1944 3085 1978
rect 3123 1944 3157 1978
rect 3195 1944 3229 1978
rect 3051 1870 3085 1904
rect 3123 1870 3157 1904
rect 3195 1870 3229 1904
rect 3051 1796 3085 1830
rect 3123 1796 3157 1830
rect 3195 1796 3229 1830
rect 3051 1722 3085 1756
rect 3123 1722 3157 1756
rect 3195 1722 3229 1756
rect 3051 1648 3085 1682
rect 3123 1648 3157 1682
rect 3195 1648 3229 1682
rect 3051 1574 3085 1608
rect 3123 1574 3157 1608
rect 3195 1574 3229 1608
rect 2872 1144 2978 1250
rect 3619 4092 3653 4118
rect 3547 4082 3725 4092
rect 3547 4048 3551 4082
rect 3551 4048 3619 4082
rect 3619 4048 3653 4082
rect 3653 4048 3721 4082
rect 3721 4048 3725 4082
rect 3547 4014 3725 4048
rect 3547 3980 3551 4014
rect 3551 3980 3619 4014
rect 3619 3980 3653 4014
rect 3653 3980 3721 4014
rect 3721 3980 3725 4014
rect 3547 3946 3725 3980
rect 3547 3912 3551 3946
rect 3551 3912 3619 3946
rect 3619 3912 3653 3946
rect 3653 3912 3721 3946
rect 3721 3912 3725 3946
rect 3547 3878 3725 3912
rect 3547 3844 3551 3878
rect 3551 3844 3619 3878
rect 3619 3844 3653 3878
rect 3653 3844 3721 3878
rect 3721 3844 3725 3878
rect 3547 3810 3725 3844
rect 3547 3776 3551 3810
rect 3551 3776 3619 3810
rect 3619 3776 3653 3810
rect 3653 3776 3721 3810
rect 3721 3776 3725 3810
rect 3547 3742 3725 3776
rect 3547 3708 3551 3742
rect 3551 3708 3619 3742
rect 3619 3708 3653 3742
rect 3653 3708 3721 3742
rect 3721 3708 3725 3742
rect 3547 3674 3725 3708
rect 3547 3640 3551 3674
rect 3551 3640 3619 3674
rect 3619 3640 3653 3674
rect 3653 3640 3721 3674
rect 3721 3640 3725 3674
rect 3547 3606 3725 3640
rect 3547 3572 3551 3606
rect 3551 3572 3619 3606
rect 3619 3572 3653 3606
rect 3653 3572 3721 3606
rect 3721 3572 3725 3606
rect 3547 3538 3725 3572
rect 3547 3504 3551 3538
rect 3551 3504 3619 3538
rect 3619 3504 3653 3538
rect 3653 3504 3721 3538
rect 3721 3504 3725 3538
rect 3547 3470 3725 3504
rect 3547 3436 3551 3470
rect 3551 3436 3619 3470
rect 3619 3436 3653 3470
rect 3653 3436 3721 3470
rect 3721 3436 3725 3470
rect 3547 3402 3725 3436
rect 3547 3368 3551 3402
rect 3551 3368 3619 3402
rect 3619 3368 3653 3402
rect 3653 3368 3721 3402
rect 3721 3368 3725 3402
rect 3547 3334 3725 3368
rect 3547 3300 3551 3334
rect 3551 3300 3619 3334
rect 3619 3300 3653 3334
rect 3653 3300 3721 3334
rect 3721 3300 3725 3334
rect 3547 3266 3725 3300
rect 3547 3232 3551 3266
rect 3551 3232 3619 3266
rect 3619 3232 3653 3266
rect 3653 3232 3721 3266
rect 3721 3232 3725 3266
rect 3547 3198 3725 3232
rect 3547 3194 3551 3198
rect 3551 3194 3619 3198
rect 3619 3194 3653 3198
rect 3653 3194 3721 3198
rect 3721 3194 3725 3198
rect 3619 3164 3653 3182
rect 3619 3148 3653 3164
rect 3547 3074 3581 3108
rect 3619 3074 3653 3108
rect 3691 3074 3725 3108
rect 3547 2994 3581 3028
rect 3619 2994 3653 3028
rect 3691 2994 3725 3028
rect 3547 2914 3581 2948
rect 3619 2914 3653 2948
rect 3691 2914 3725 2948
rect 3547 2834 3581 2868
rect 3619 2834 3653 2868
rect 3691 2834 3725 2868
rect 3547 2754 3581 2788
rect 3619 2754 3653 2788
rect 3691 2754 3725 2788
rect 3547 2674 3581 2708
rect 3619 2674 3653 2708
rect 3691 2674 3725 2708
rect 3547 2594 3581 2628
rect 3619 2594 3653 2628
rect 3691 2594 3725 2628
rect 3619 2540 3653 2556
rect 3619 2522 3653 2540
rect 3547 2506 3551 2518
rect 3551 2506 3619 2518
rect 3619 2506 3653 2518
rect 3653 2506 3721 2518
rect 3721 2506 3725 2518
rect 3547 2472 3725 2506
rect 3547 2438 3551 2472
rect 3551 2438 3619 2472
rect 3619 2438 3653 2472
rect 3653 2438 3721 2472
rect 3721 2438 3725 2472
rect 3547 2404 3725 2438
rect 3547 2370 3551 2404
rect 3551 2370 3619 2404
rect 3619 2370 3653 2404
rect 3653 2370 3721 2404
rect 3721 2370 3725 2404
rect 3547 2336 3725 2370
rect 3547 2302 3551 2336
rect 3551 2302 3619 2336
rect 3619 2302 3653 2336
rect 3653 2302 3721 2336
rect 3721 2302 3725 2336
rect 3547 2268 3725 2302
rect 3547 2234 3551 2268
rect 3551 2234 3619 2268
rect 3619 2234 3653 2268
rect 3653 2234 3721 2268
rect 3721 2234 3725 2268
rect 3547 2200 3725 2234
rect 3547 2166 3551 2200
rect 3551 2166 3619 2200
rect 3619 2166 3653 2200
rect 3653 2166 3721 2200
rect 3721 2166 3725 2200
rect 3547 2132 3725 2166
rect 3547 2098 3551 2132
rect 3551 2098 3619 2132
rect 3619 2098 3653 2132
rect 3653 2098 3721 2132
rect 3721 2098 3725 2132
rect 3547 2064 3725 2098
rect 3547 2030 3551 2064
rect 3551 2030 3619 2064
rect 3619 2030 3653 2064
rect 3653 2030 3721 2064
rect 3721 2030 3725 2064
rect 3547 1996 3725 2030
rect 3547 1962 3551 1996
rect 3551 1962 3619 1996
rect 3619 1962 3653 1996
rect 3653 1962 3721 1996
rect 3721 1962 3725 1996
rect 3547 1928 3725 1962
rect 3547 1894 3551 1928
rect 3551 1894 3619 1928
rect 3619 1894 3653 1928
rect 3653 1894 3721 1928
rect 3721 1894 3725 1928
rect 3547 1860 3725 1894
rect 3547 1826 3551 1860
rect 3551 1826 3619 1860
rect 3619 1826 3653 1860
rect 3653 1826 3721 1860
rect 3721 1826 3725 1860
rect 3547 1792 3725 1826
rect 3547 1758 3551 1792
rect 3551 1758 3619 1792
rect 3619 1758 3653 1792
rect 3653 1758 3721 1792
rect 3721 1758 3725 1792
rect 3547 1724 3725 1758
rect 3547 1690 3551 1724
rect 3551 1690 3619 1724
rect 3619 1690 3653 1724
rect 3653 1690 3721 1724
rect 3721 1690 3725 1724
rect 3547 1656 3725 1690
rect 3547 1622 3551 1656
rect 3551 1622 3619 1656
rect 3619 1622 3653 1656
rect 3653 1622 3721 1656
rect 3721 1622 3725 1656
rect 3547 1620 3725 1622
rect 3619 1586 3653 1620
rect 3302 1144 3408 1250
rect 4043 4064 4077 4098
rect 4115 4064 4149 4098
rect 4187 4064 4221 4098
rect 4043 3991 4077 4025
rect 4115 3991 4149 4025
rect 4187 3991 4221 4025
rect 4043 3918 4077 3952
rect 4115 3918 4149 3952
rect 4187 3918 4221 3952
rect 4043 3845 4077 3879
rect 4115 3845 4149 3879
rect 4187 3845 4221 3879
rect 4043 3772 4077 3806
rect 4115 3772 4149 3806
rect 4187 3772 4221 3806
rect 4043 3699 4077 3733
rect 4115 3699 4149 3733
rect 4187 3699 4221 3733
rect 4043 3626 4077 3660
rect 4115 3626 4149 3660
rect 4187 3626 4221 3660
rect 4043 3553 4077 3587
rect 4115 3553 4149 3587
rect 4187 3553 4221 3587
rect 4043 3480 4077 3514
rect 4115 3480 4149 3514
rect 4187 3480 4221 3514
rect 4043 3407 4077 3441
rect 4115 3407 4149 3441
rect 4187 3407 4221 3441
rect 4043 3334 4077 3368
rect 4115 3334 4149 3368
rect 4187 3334 4221 3368
rect 4043 3261 4077 3295
rect 4115 3261 4149 3295
rect 4187 3261 4221 3295
rect 4043 3188 4077 3222
rect 4115 3188 4149 3222
rect 4187 3188 4221 3222
rect 4043 3115 4077 3149
rect 4115 3115 4149 3149
rect 4187 3115 4221 3149
rect 4043 3042 4077 3076
rect 4115 3042 4149 3076
rect 4187 3042 4221 3076
rect 4043 2969 4077 3003
rect 4115 2969 4149 3003
rect 4187 2969 4221 3003
rect 4043 2896 4077 2930
rect 4115 2896 4149 2930
rect 4187 2896 4221 2930
rect 4043 2823 4077 2857
rect 4115 2823 4149 2857
rect 4187 2823 4221 2857
rect 4043 2750 4077 2784
rect 4115 2750 4149 2784
rect 4187 2750 4221 2784
rect 4043 2677 4077 2711
rect 4115 2677 4149 2711
rect 4187 2677 4221 2711
rect 4043 2604 4077 2638
rect 4115 2604 4149 2638
rect 4187 2604 4221 2638
rect 4043 2531 4077 2565
rect 4115 2531 4149 2565
rect 4187 2531 4221 2565
rect 4043 2458 4077 2492
rect 4115 2458 4149 2492
rect 4187 2458 4221 2492
rect 4043 2385 4077 2419
rect 4115 2385 4149 2419
rect 4187 2385 4221 2419
rect 4043 2312 4077 2346
rect 4115 2312 4149 2346
rect 4187 2312 4221 2346
rect 4043 2239 4077 2273
rect 4115 2239 4149 2273
rect 4187 2239 4221 2273
rect 4043 2166 4077 2200
rect 4115 2166 4149 2200
rect 4187 2166 4221 2200
rect 4043 2092 4077 2126
rect 4115 2092 4149 2126
rect 4187 2092 4221 2126
rect 4043 2018 4077 2052
rect 4115 2018 4149 2052
rect 4187 2018 4221 2052
rect 4043 1944 4077 1978
rect 4115 1944 4149 1978
rect 4187 1944 4221 1978
rect 4043 1870 4077 1904
rect 4115 1870 4149 1904
rect 4187 1870 4221 1904
rect 4043 1796 4077 1830
rect 4115 1796 4149 1830
rect 4187 1796 4221 1830
rect 4043 1722 4077 1756
rect 4115 1722 4149 1756
rect 4187 1722 4221 1756
rect 4043 1648 4077 1682
rect 4115 1648 4149 1682
rect 4187 1648 4221 1682
rect 4043 1574 4077 1608
rect 4115 1574 4149 1608
rect 4187 1574 4221 1608
rect 3864 1144 3970 1250
rect 4611 4092 4645 4118
rect 4539 4082 4717 4092
rect 4539 4048 4543 4082
rect 4543 4048 4611 4082
rect 4611 4048 4645 4082
rect 4645 4048 4713 4082
rect 4713 4048 4717 4082
rect 4539 4014 4717 4048
rect 4539 3980 4543 4014
rect 4543 3980 4611 4014
rect 4611 3980 4645 4014
rect 4645 3980 4713 4014
rect 4713 3980 4717 4014
rect 4539 3946 4717 3980
rect 4539 3912 4543 3946
rect 4543 3912 4611 3946
rect 4611 3912 4645 3946
rect 4645 3912 4713 3946
rect 4713 3912 4717 3946
rect 4539 3878 4717 3912
rect 4539 3844 4543 3878
rect 4543 3844 4611 3878
rect 4611 3844 4645 3878
rect 4645 3844 4713 3878
rect 4713 3844 4717 3878
rect 4539 3810 4717 3844
rect 4539 3776 4543 3810
rect 4543 3776 4611 3810
rect 4611 3776 4645 3810
rect 4645 3776 4713 3810
rect 4713 3776 4717 3810
rect 4539 3742 4717 3776
rect 4539 3708 4543 3742
rect 4543 3708 4611 3742
rect 4611 3708 4645 3742
rect 4645 3708 4713 3742
rect 4713 3708 4717 3742
rect 4539 3674 4717 3708
rect 4539 3640 4543 3674
rect 4543 3640 4611 3674
rect 4611 3640 4645 3674
rect 4645 3640 4713 3674
rect 4713 3640 4717 3674
rect 4539 3606 4717 3640
rect 4539 3572 4543 3606
rect 4543 3572 4611 3606
rect 4611 3572 4645 3606
rect 4645 3572 4713 3606
rect 4713 3572 4717 3606
rect 4539 3538 4717 3572
rect 4539 3504 4543 3538
rect 4543 3504 4611 3538
rect 4611 3504 4645 3538
rect 4645 3504 4713 3538
rect 4713 3504 4717 3538
rect 4539 3470 4717 3504
rect 4539 3436 4543 3470
rect 4543 3436 4611 3470
rect 4611 3436 4645 3470
rect 4645 3436 4713 3470
rect 4713 3436 4717 3470
rect 4539 3402 4717 3436
rect 4539 3368 4543 3402
rect 4543 3368 4611 3402
rect 4611 3368 4645 3402
rect 4645 3368 4713 3402
rect 4713 3368 4717 3402
rect 4539 3334 4717 3368
rect 4539 3300 4543 3334
rect 4543 3300 4611 3334
rect 4611 3300 4645 3334
rect 4645 3300 4713 3334
rect 4713 3300 4717 3334
rect 4539 3266 4717 3300
rect 4539 3232 4543 3266
rect 4543 3232 4611 3266
rect 4611 3232 4645 3266
rect 4645 3232 4713 3266
rect 4713 3232 4717 3266
rect 4539 3198 4717 3232
rect 4539 3194 4543 3198
rect 4543 3194 4611 3198
rect 4611 3194 4645 3198
rect 4645 3194 4713 3198
rect 4713 3194 4717 3198
rect 4611 3164 4645 3182
rect 4611 3148 4645 3164
rect 4539 3074 4573 3108
rect 4611 3074 4645 3108
rect 4683 3074 4717 3108
rect 4539 2994 4573 3028
rect 4611 2994 4645 3028
rect 4683 2994 4717 3028
rect 4539 2914 4573 2948
rect 4611 2914 4645 2948
rect 4683 2914 4717 2948
rect 4539 2834 4573 2868
rect 4611 2834 4645 2868
rect 4683 2834 4717 2868
rect 4539 2754 4573 2788
rect 4611 2754 4645 2788
rect 4683 2754 4717 2788
rect 4539 2674 4573 2708
rect 4611 2674 4645 2708
rect 4683 2674 4717 2708
rect 4539 2594 4573 2628
rect 4611 2594 4645 2628
rect 4683 2594 4717 2628
rect 4611 2540 4645 2556
rect 4611 2522 4645 2540
rect 4539 2506 4543 2518
rect 4543 2506 4611 2518
rect 4611 2506 4645 2518
rect 4645 2506 4713 2518
rect 4713 2506 4717 2518
rect 4539 2472 4717 2506
rect 4539 2438 4543 2472
rect 4543 2438 4611 2472
rect 4611 2438 4645 2472
rect 4645 2438 4713 2472
rect 4713 2438 4717 2472
rect 4539 2404 4717 2438
rect 4539 2370 4543 2404
rect 4543 2370 4611 2404
rect 4611 2370 4645 2404
rect 4645 2370 4713 2404
rect 4713 2370 4717 2404
rect 4539 2336 4717 2370
rect 4539 2302 4543 2336
rect 4543 2302 4611 2336
rect 4611 2302 4645 2336
rect 4645 2302 4713 2336
rect 4713 2302 4717 2336
rect 4539 2268 4717 2302
rect 4539 2234 4543 2268
rect 4543 2234 4611 2268
rect 4611 2234 4645 2268
rect 4645 2234 4713 2268
rect 4713 2234 4717 2268
rect 4539 2200 4717 2234
rect 4539 2166 4543 2200
rect 4543 2166 4611 2200
rect 4611 2166 4645 2200
rect 4645 2166 4713 2200
rect 4713 2166 4717 2200
rect 4539 2132 4717 2166
rect 4539 2098 4543 2132
rect 4543 2098 4611 2132
rect 4611 2098 4645 2132
rect 4645 2098 4713 2132
rect 4713 2098 4717 2132
rect 4539 2064 4717 2098
rect 4539 2030 4543 2064
rect 4543 2030 4611 2064
rect 4611 2030 4645 2064
rect 4645 2030 4713 2064
rect 4713 2030 4717 2064
rect 4539 1996 4717 2030
rect 4539 1962 4543 1996
rect 4543 1962 4611 1996
rect 4611 1962 4645 1996
rect 4645 1962 4713 1996
rect 4713 1962 4717 1996
rect 4539 1928 4717 1962
rect 4539 1894 4543 1928
rect 4543 1894 4611 1928
rect 4611 1894 4645 1928
rect 4645 1894 4713 1928
rect 4713 1894 4717 1928
rect 4539 1860 4717 1894
rect 4539 1826 4543 1860
rect 4543 1826 4611 1860
rect 4611 1826 4645 1860
rect 4645 1826 4713 1860
rect 4713 1826 4717 1860
rect 4539 1792 4717 1826
rect 4539 1758 4543 1792
rect 4543 1758 4611 1792
rect 4611 1758 4645 1792
rect 4645 1758 4713 1792
rect 4713 1758 4717 1792
rect 4539 1724 4717 1758
rect 4539 1690 4543 1724
rect 4543 1690 4611 1724
rect 4611 1690 4645 1724
rect 4645 1690 4713 1724
rect 4713 1690 4717 1724
rect 4539 1656 4717 1690
rect 4539 1622 4543 1656
rect 4543 1622 4611 1656
rect 4611 1622 4645 1656
rect 4645 1622 4713 1656
rect 4713 1622 4717 1656
rect 4539 1620 4717 1622
rect 4611 1586 4645 1620
rect 4294 1144 4400 1250
rect 5035 4064 5069 4098
rect 5107 4064 5141 4098
rect 5179 4064 5213 4098
rect 5035 3991 5069 4025
rect 5107 3991 5141 4025
rect 5179 3991 5213 4025
rect 5035 3918 5069 3952
rect 5107 3918 5141 3952
rect 5179 3918 5213 3952
rect 5035 3845 5069 3879
rect 5107 3845 5141 3879
rect 5179 3845 5213 3879
rect 5035 3772 5069 3806
rect 5107 3772 5141 3806
rect 5179 3772 5213 3806
rect 5035 3699 5069 3733
rect 5107 3699 5141 3733
rect 5179 3699 5213 3733
rect 5035 3626 5069 3660
rect 5107 3626 5141 3660
rect 5179 3626 5213 3660
rect 5035 3553 5069 3587
rect 5107 3553 5141 3587
rect 5179 3553 5213 3587
rect 5035 3480 5069 3514
rect 5107 3480 5141 3514
rect 5179 3480 5213 3514
rect 5035 3407 5069 3441
rect 5107 3407 5141 3441
rect 5179 3407 5213 3441
rect 5035 3334 5069 3368
rect 5107 3334 5141 3368
rect 5179 3334 5213 3368
rect 5035 3261 5069 3295
rect 5107 3261 5141 3295
rect 5179 3261 5213 3295
rect 5035 3188 5069 3222
rect 5107 3188 5141 3222
rect 5179 3188 5213 3222
rect 5035 3115 5069 3149
rect 5107 3115 5141 3149
rect 5179 3115 5213 3149
rect 5035 3042 5069 3076
rect 5107 3042 5141 3076
rect 5179 3042 5213 3076
rect 5035 2969 5069 3003
rect 5107 2969 5141 3003
rect 5179 2969 5213 3003
rect 5035 2896 5069 2930
rect 5107 2896 5141 2930
rect 5179 2896 5213 2930
rect 5035 2823 5069 2857
rect 5107 2823 5141 2857
rect 5179 2823 5213 2857
rect 5035 2750 5069 2784
rect 5107 2750 5141 2784
rect 5179 2750 5213 2784
rect 5035 2677 5069 2711
rect 5107 2677 5141 2711
rect 5179 2677 5213 2711
rect 5035 2604 5069 2638
rect 5107 2604 5141 2638
rect 5179 2604 5213 2638
rect 5035 2531 5069 2565
rect 5107 2531 5141 2565
rect 5179 2531 5213 2565
rect 5035 2458 5069 2492
rect 5107 2458 5141 2492
rect 5179 2458 5213 2492
rect 5035 2385 5069 2419
rect 5107 2385 5141 2419
rect 5179 2385 5213 2419
rect 5035 2312 5069 2346
rect 5107 2312 5141 2346
rect 5179 2312 5213 2346
rect 5035 2239 5069 2273
rect 5107 2239 5141 2273
rect 5179 2239 5213 2273
rect 5035 2166 5069 2200
rect 5107 2166 5141 2200
rect 5179 2166 5213 2200
rect 5035 2092 5069 2126
rect 5107 2092 5141 2126
rect 5179 2092 5213 2126
rect 5035 2018 5069 2052
rect 5107 2018 5141 2052
rect 5179 2018 5213 2052
rect 5035 1944 5069 1978
rect 5107 1944 5141 1978
rect 5179 1944 5213 1978
rect 5035 1870 5069 1904
rect 5107 1870 5141 1904
rect 5179 1870 5213 1904
rect 5035 1796 5069 1830
rect 5107 1796 5141 1830
rect 5179 1796 5213 1830
rect 5035 1722 5069 1756
rect 5107 1722 5141 1756
rect 5179 1722 5213 1756
rect 5035 1648 5069 1682
rect 5107 1648 5141 1682
rect 5179 1648 5213 1682
rect 5035 1574 5069 1608
rect 5107 1574 5141 1608
rect 5179 1574 5213 1608
rect 4856 1144 4962 1250
rect 5603 4092 5637 4118
rect 5531 4082 5709 4092
rect 5531 4048 5535 4082
rect 5535 4048 5603 4082
rect 5603 4048 5637 4082
rect 5637 4048 5705 4082
rect 5705 4048 5709 4082
rect 5531 4014 5709 4048
rect 5531 3980 5535 4014
rect 5535 3980 5603 4014
rect 5603 3980 5637 4014
rect 5637 3980 5705 4014
rect 5705 3980 5709 4014
rect 5531 3946 5709 3980
rect 5531 3912 5535 3946
rect 5535 3912 5603 3946
rect 5603 3912 5637 3946
rect 5637 3912 5705 3946
rect 5705 3912 5709 3946
rect 5531 3878 5709 3912
rect 5531 3844 5535 3878
rect 5535 3844 5603 3878
rect 5603 3844 5637 3878
rect 5637 3844 5705 3878
rect 5705 3844 5709 3878
rect 5531 3810 5709 3844
rect 5531 3776 5535 3810
rect 5535 3776 5603 3810
rect 5603 3776 5637 3810
rect 5637 3776 5705 3810
rect 5705 3776 5709 3810
rect 5531 3742 5709 3776
rect 5531 3708 5535 3742
rect 5535 3708 5603 3742
rect 5603 3708 5637 3742
rect 5637 3708 5705 3742
rect 5705 3708 5709 3742
rect 5531 3674 5709 3708
rect 5531 3640 5535 3674
rect 5535 3640 5603 3674
rect 5603 3640 5637 3674
rect 5637 3640 5705 3674
rect 5705 3640 5709 3674
rect 5531 3606 5709 3640
rect 5531 3572 5535 3606
rect 5535 3572 5603 3606
rect 5603 3572 5637 3606
rect 5637 3572 5705 3606
rect 5705 3572 5709 3606
rect 5531 3538 5709 3572
rect 5531 3504 5535 3538
rect 5535 3504 5603 3538
rect 5603 3504 5637 3538
rect 5637 3504 5705 3538
rect 5705 3504 5709 3538
rect 5531 3470 5709 3504
rect 5531 3436 5535 3470
rect 5535 3436 5603 3470
rect 5603 3436 5637 3470
rect 5637 3436 5705 3470
rect 5705 3436 5709 3470
rect 5531 3402 5709 3436
rect 5531 3368 5535 3402
rect 5535 3368 5603 3402
rect 5603 3368 5637 3402
rect 5637 3368 5705 3402
rect 5705 3368 5709 3402
rect 5531 3334 5709 3368
rect 5531 3300 5535 3334
rect 5535 3300 5603 3334
rect 5603 3300 5637 3334
rect 5637 3300 5705 3334
rect 5705 3300 5709 3334
rect 5531 3266 5709 3300
rect 5531 3232 5535 3266
rect 5535 3232 5603 3266
rect 5603 3232 5637 3266
rect 5637 3232 5705 3266
rect 5705 3232 5709 3266
rect 5531 3198 5709 3232
rect 5531 3194 5535 3198
rect 5535 3194 5603 3198
rect 5603 3194 5637 3198
rect 5637 3194 5705 3198
rect 5705 3194 5709 3198
rect 5603 3164 5637 3182
rect 5603 3148 5637 3164
rect 5531 3074 5565 3108
rect 5603 3074 5637 3108
rect 5675 3074 5709 3108
rect 5531 2994 5565 3028
rect 5603 2994 5637 3028
rect 5675 2994 5709 3028
rect 5531 2914 5565 2948
rect 5603 2914 5637 2948
rect 5675 2914 5709 2948
rect 5531 2834 5565 2868
rect 5603 2834 5637 2868
rect 5675 2834 5709 2868
rect 5531 2754 5565 2788
rect 5603 2754 5637 2788
rect 5675 2754 5709 2788
rect 5531 2674 5565 2708
rect 5603 2674 5637 2708
rect 5675 2674 5709 2708
rect 5531 2594 5565 2628
rect 5603 2594 5637 2628
rect 5675 2594 5709 2628
rect 5603 2540 5637 2556
rect 5603 2522 5637 2540
rect 5531 2506 5535 2518
rect 5535 2506 5603 2518
rect 5603 2506 5637 2518
rect 5637 2506 5705 2518
rect 5705 2506 5709 2518
rect 5531 2472 5709 2506
rect 5531 2438 5535 2472
rect 5535 2438 5603 2472
rect 5603 2438 5637 2472
rect 5637 2438 5705 2472
rect 5705 2438 5709 2472
rect 5531 2404 5709 2438
rect 5531 2370 5535 2404
rect 5535 2370 5603 2404
rect 5603 2370 5637 2404
rect 5637 2370 5705 2404
rect 5705 2370 5709 2404
rect 5531 2336 5709 2370
rect 5531 2302 5535 2336
rect 5535 2302 5603 2336
rect 5603 2302 5637 2336
rect 5637 2302 5705 2336
rect 5705 2302 5709 2336
rect 5531 2268 5709 2302
rect 5531 2234 5535 2268
rect 5535 2234 5603 2268
rect 5603 2234 5637 2268
rect 5637 2234 5705 2268
rect 5705 2234 5709 2268
rect 5531 2200 5709 2234
rect 5531 2166 5535 2200
rect 5535 2166 5603 2200
rect 5603 2166 5637 2200
rect 5637 2166 5705 2200
rect 5705 2166 5709 2200
rect 5531 2132 5709 2166
rect 5531 2098 5535 2132
rect 5535 2098 5603 2132
rect 5603 2098 5637 2132
rect 5637 2098 5705 2132
rect 5705 2098 5709 2132
rect 5531 2064 5709 2098
rect 5531 2030 5535 2064
rect 5535 2030 5603 2064
rect 5603 2030 5637 2064
rect 5637 2030 5705 2064
rect 5705 2030 5709 2064
rect 5531 1996 5709 2030
rect 5531 1962 5535 1996
rect 5535 1962 5603 1996
rect 5603 1962 5637 1996
rect 5637 1962 5705 1996
rect 5705 1962 5709 1996
rect 5531 1928 5709 1962
rect 5531 1894 5535 1928
rect 5535 1894 5603 1928
rect 5603 1894 5637 1928
rect 5637 1894 5705 1928
rect 5705 1894 5709 1928
rect 5531 1860 5709 1894
rect 5531 1826 5535 1860
rect 5535 1826 5603 1860
rect 5603 1826 5637 1860
rect 5637 1826 5705 1860
rect 5705 1826 5709 1860
rect 5531 1792 5709 1826
rect 5531 1758 5535 1792
rect 5535 1758 5603 1792
rect 5603 1758 5637 1792
rect 5637 1758 5705 1792
rect 5705 1758 5709 1792
rect 5531 1724 5709 1758
rect 5531 1690 5535 1724
rect 5535 1690 5603 1724
rect 5603 1690 5637 1724
rect 5637 1690 5705 1724
rect 5705 1690 5709 1724
rect 5531 1656 5709 1690
rect 5531 1622 5535 1656
rect 5535 1622 5603 1656
rect 5603 1622 5637 1656
rect 5637 1622 5705 1656
rect 5705 1622 5709 1656
rect 5531 1620 5709 1622
rect 5603 1586 5637 1620
rect 5286 1144 5392 1250
rect 6027 4064 6061 4098
rect 6099 4064 6133 4098
rect 6171 4064 6205 4098
rect 6027 3991 6061 4025
rect 6099 3991 6133 4025
rect 6171 3991 6205 4025
rect 6027 3918 6061 3952
rect 6099 3918 6133 3952
rect 6171 3918 6205 3952
rect 6027 3845 6061 3879
rect 6099 3845 6133 3879
rect 6171 3845 6205 3879
rect 6027 3772 6061 3806
rect 6099 3772 6133 3806
rect 6171 3772 6205 3806
rect 6027 3699 6061 3733
rect 6099 3699 6133 3733
rect 6171 3699 6205 3733
rect 6027 3626 6061 3660
rect 6099 3626 6133 3660
rect 6171 3626 6205 3660
rect 6027 3553 6061 3587
rect 6099 3553 6133 3587
rect 6171 3553 6205 3587
rect 6027 3480 6061 3514
rect 6099 3480 6133 3514
rect 6171 3480 6205 3514
rect 6027 3407 6061 3441
rect 6099 3407 6133 3441
rect 6171 3407 6205 3441
rect 6027 3334 6061 3368
rect 6099 3334 6133 3368
rect 6171 3334 6205 3368
rect 6027 3261 6061 3295
rect 6099 3261 6133 3295
rect 6171 3261 6205 3295
rect 6027 3188 6061 3222
rect 6099 3188 6133 3222
rect 6171 3188 6205 3222
rect 6027 3115 6061 3149
rect 6099 3115 6133 3149
rect 6171 3115 6205 3149
rect 6027 3042 6061 3076
rect 6099 3042 6133 3076
rect 6171 3042 6205 3076
rect 6027 2969 6061 3003
rect 6099 2969 6133 3003
rect 6171 2969 6205 3003
rect 6027 2896 6061 2930
rect 6099 2896 6133 2930
rect 6171 2896 6205 2930
rect 6027 2823 6061 2857
rect 6099 2823 6133 2857
rect 6171 2823 6205 2857
rect 6027 2750 6061 2784
rect 6099 2750 6133 2784
rect 6171 2750 6205 2784
rect 6027 2677 6061 2711
rect 6099 2677 6133 2711
rect 6171 2677 6205 2711
rect 6027 2604 6061 2638
rect 6099 2604 6133 2638
rect 6171 2604 6205 2638
rect 6027 2531 6061 2565
rect 6099 2531 6133 2565
rect 6171 2531 6205 2565
rect 6027 2458 6061 2492
rect 6099 2458 6133 2492
rect 6171 2458 6205 2492
rect 6027 2385 6061 2419
rect 6099 2385 6133 2419
rect 6171 2385 6205 2419
rect 6027 2312 6061 2346
rect 6099 2312 6133 2346
rect 6171 2312 6205 2346
rect 6027 2239 6061 2273
rect 6099 2239 6133 2273
rect 6171 2239 6205 2273
rect 6027 2166 6061 2200
rect 6099 2166 6133 2200
rect 6171 2166 6205 2200
rect 6027 2092 6061 2126
rect 6099 2092 6133 2126
rect 6171 2092 6205 2126
rect 6027 2018 6061 2052
rect 6099 2018 6133 2052
rect 6171 2018 6205 2052
rect 6027 1944 6061 1978
rect 6099 1944 6133 1978
rect 6171 1944 6205 1978
rect 6027 1870 6061 1904
rect 6099 1870 6133 1904
rect 6171 1870 6205 1904
rect 6027 1796 6061 1830
rect 6099 1796 6133 1830
rect 6171 1796 6205 1830
rect 6027 1722 6061 1756
rect 6099 1722 6133 1756
rect 6171 1722 6205 1756
rect 6027 1648 6061 1682
rect 6099 1648 6133 1682
rect 6171 1648 6205 1682
rect 6027 1574 6061 1608
rect 6099 1574 6133 1608
rect 6171 1574 6205 1608
rect 5848 1144 5954 1250
rect 6595 4092 6629 4118
rect 6523 4082 6701 4092
rect 6523 4048 6527 4082
rect 6527 4048 6595 4082
rect 6595 4048 6629 4082
rect 6629 4048 6697 4082
rect 6697 4048 6701 4082
rect 6523 4014 6701 4048
rect 6523 3980 6527 4014
rect 6527 3980 6595 4014
rect 6595 3980 6629 4014
rect 6629 3980 6697 4014
rect 6697 3980 6701 4014
rect 6523 3946 6701 3980
rect 6523 3912 6527 3946
rect 6527 3912 6595 3946
rect 6595 3912 6629 3946
rect 6629 3912 6697 3946
rect 6697 3912 6701 3946
rect 6523 3878 6701 3912
rect 6523 3844 6527 3878
rect 6527 3844 6595 3878
rect 6595 3844 6629 3878
rect 6629 3844 6697 3878
rect 6697 3844 6701 3878
rect 6523 3810 6701 3844
rect 6523 3776 6527 3810
rect 6527 3776 6595 3810
rect 6595 3776 6629 3810
rect 6629 3776 6697 3810
rect 6697 3776 6701 3810
rect 6523 3742 6701 3776
rect 6523 3708 6527 3742
rect 6527 3708 6595 3742
rect 6595 3708 6629 3742
rect 6629 3708 6697 3742
rect 6697 3708 6701 3742
rect 6523 3674 6701 3708
rect 6523 3640 6527 3674
rect 6527 3640 6595 3674
rect 6595 3640 6629 3674
rect 6629 3640 6697 3674
rect 6697 3640 6701 3674
rect 6523 3606 6701 3640
rect 6523 3572 6527 3606
rect 6527 3572 6595 3606
rect 6595 3572 6629 3606
rect 6629 3572 6697 3606
rect 6697 3572 6701 3606
rect 6523 3538 6701 3572
rect 6523 3504 6527 3538
rect 6527 3504 6595 3538
rect 6595 3504 6629 3538
rect 6629 3504 6697 3538
rect 6697 3504 6701 3538
rect 6523 3470 6701 3504
rect 6523 3436 6527 3470
rect 6527 3436 6595 3470
rect 6595 3436 6629 3470
rect 6629 3436 6697 3470
rect 6697 3436 6701 3470
rect 6523 3402 6701 3436
rect 6523 3368 6527 3402
rect 6527 3368 6595 3402
rect 6595 3368 6629 3402
rect 6629 3368 6697 3402
rect 6697 3368 6701 3402
rect 6523 3334 6701 3368
rect 6523 3300 6527 3334
rect 6527 3300 6595 3334
rect 6595 3300 6629 3334
rect 6629 3300 6697 3334
rect 6697 3300 6701 3334
rect 6523 3266 6701 3300
rect 6523 3232 6527 3266
rect 6527 3232 6595 3266
rect 6595 3232 6629 3266
rect 6629 3232 6697 3266
rect 6697 3232 6701 3266
rect 6523 3198 6701 3232
rect 6523 3194 6527 3198
rect 6527 3194 6595 3198
rect 6595 3194 6629 3198
rect 6629 3194 6697 3198
rect 6697 3194 6701 3198
rect 6595 3164 6629 3182
rect 6595 3148 6629 3164
rect 6523 3074 6557 3108
rect 6595 3074 6629 3108
rect 6667 3074 6701 3108
rect 6523 2994 6557 3028
rect 6595 2994 6629 3028
rect 6667 2994 6701 3028
rect 6523 2914 6557 2948
rect 6595 2914 6629 2948
rect 6667 2914 6701 2948
rect 6523 2834 6557 2868
rect 6595 2834 6629 2868
rect 6667 2834 6701 2868
rect 6523 2754 6557 2788
rect 6595 2754 6629 2788
rect 6667 2754 6701 2788
rect 6523 2674 6557 2708
rect 6595 2674 6629 2708
rect 6667 2674 6701 2708
rect 6523 2594 6557 2628
rect 6595 2594 6629 2628
rect 6667 2594 6701 2628
rect 6595 2540 6629 2556
rect 6595 2522 6629 2540
rect 6523 2506 6527 2518
rect 6527 2506 6595 2518
rect 6595 2506 6629 2518
rect 6629 2506 6697 2518
rect 6697 2506 6701 2518
rect 6523 2472 6701 2506
rect 6523 2438 6527 2472
rect 6527 2438 6595 2472
rect 6595 2438 6629 2472
rect 6629 2438 6697 2472
rect 6697 2438 6701 2472
rect 6523 2404 6701 2438
rect 6523 2370 6527 2404
rect 6527 2370 6595 2404
rect 6595 2370 6629 2404
rect 6629 2370 6697 2404
rect 6697 2370 6701 2404
rect 6523 2336 6701 2370
rect 6523 2302 6527 2336
rect 6527 2302 6595 2336
rect 6595 2302 6629 2336
rect 6629 2302 6697 2336
rect 6697 2302 6701 2336
rect 6523 2268 6701 2302
rect 6523 2234 6527 2268
rect 6527 2234 6595 2268
rect 6595 2234 6629 2268
rect 6629 2234 6697 2268
rect 6697 2234 6701 2268
rect 6523 2200 6701 2234
rect 6523 2166 6527 2200
rect 6527 2166 6595 2200
rect 6595 2166 6629 2200
rect 6629 2166 6697 2200
rect 6697 2166 6701 2200
rect 6523 2132 6701 2166
rect 6523 2098 6527 2132
rect 6527 2098 6595 2132
rect 6595 2098 6629 2132
rect 6629 2098 6697 2132
rect 6697 2098 6701 2132
rect 6523 2064 6701 2098
rect 6523 2030 6527 2064
rect 6527 2030 6595 2064
rect 6595 2030 6629 2064
rect 6629 2030 6697 2064
rect 6697 2030 6701 2064
rect 6523 1996 6701 2030
rect 6523 1962 6527 1996
rect 6527 1962 6595 1996
rect 6595 1962 6629 1996
rect 6629 1962 6697 1996
rect 6697 1962 6701 1996
rect 6523 1928 6701 1962
rect 6523 1894 6527 1928
rect 6527 1894 6595 1928
rect 6595 1894 6629 1928
rect 6629 1894 6697 1928
rect 6697 1894 6701 1928
rect 6523 1860 6701 1894
rect 6523 1826 6527 1860
rect 6527 1826 6595 1860
rect 6595 1826 6629 1860
rect 6629 1826 6697 1860
rect 6697 1826 6701 1860
rect 6523 1792 6701 1826
rect 6523 1758 6527 1792
rect 6527 1758 6595 1792
rect 6595 1758 6629 1792
rect 6629 1758 6697 1792
rect 6697 1758 6701 1792
rect 6523 1724 6701 1758
rect 6523 1690 6527 1724
rect 6527 1690 6595 1724
rect 6595 1690 6629 1724
rect 6629 1690 6697 1724
rect 6697 1690 6701 1724
rect 6523 1656 6701 1690
rect 6523 1622 6527 1656
rect 6527 1622 6595 1656
rect 6595 1622 6629 1656
rect 6629 1622 6697 1656
rect 6697 1622 6701 1656
rect 6523 1620 6701 1622
rect 6595 1586 6629 1620
rect 6278 1144 6384 1250
rect 7019 4064 7053 4098
rect 7091 4064 7125 4098
rect 7163 4064 7197 4098
rect 7019 3991 7053 4025
rect 7091 3991 7125 4025
rect 7163 3991 7197 4025
rect 7019 3918 7053 3952
rect 7091 3918 7125 3952
rect 7163 3918 7197 3952
rect 7019 3845 7053 3879
rect 7091 3845 7125 3879
rect 7163 3845 7197 3879
rect 7019 3772 7053 3806
rect 7091 3772 7125 3806
rect 7163 3772 7197 3806
rect 7019 3699 7053 3733
rect 7091 3699 7125 3733
rect 7163 3699 7197 3733
rect 7019 3626 7053 3660
rect 7091 3626 7125 3660
rect 7163 3626 7197 3660
rect 7019 3553 7053 3587
rect 7091 3553 7125 3587
rect 7163 3553 7197 3587
rect 7019 3480 7053 3514
rect 7091 3480 7125 3514
rect 7163 3480 7197 3514
rect 7019 3407 7053 3441
rect 7091 3407 7125 3441
rect 7163 3407 7197 3441
rect 7019 3334 7053 3368
rect 7091 3334 7125 3368
rect 7163 3334 7197 3368
rect 7019 3261 7053 3295
rect 7091 3261 7125 3295
rect 7163 3261 7197 3295
rect 7019 3188 7053 3222
rect 7091 3188 7125 3222
rect 7163 3188 7197 3222
rect 7019 3115 7053 3149
rect 7091 3115 7125 3149
rect 7163 3115 7197 3149
rect 7019 3042 7053 3076
rect 7091 3042 7125 3076
rect 7163 3042 7197 3076
rect 7019 2969 7053 3003
rect 7091 2969 7125 3003
rect 7163 2969 7197 3003
rect 7019 2896 7053 2930
rect 7091 2896 7125 2930
rect 7163 2896 7197 2930
rect 7019 2823 7053 2857
rect 7091 2823 7125 2857
rect 7163 2823 7197 2857
rect 7019 2750 7053 2784
rect 7091 2750 7125 2784
rect 7163 2750 7197 2784
rect 7019 2677 7053 2711
rect 7091 2677 7125 2711
rect 7163 2677 7197 2711
rect 7019 2604 7053 2638
rect 7091 2604 7125 2638
rect 7163 2604 7197 2638
rect 7019 2531 7053 2565
rect 7091 2531 7125 2565
rect 7163 2531 7197 2565
rect 7019 2458 7053 2492
rect 7091 2458 7125 2492
rect 7163 2458 7197 2492
rect 7019 2385 7053 2419
rect 7091 2385 7125 2419
rect 7163 2385 7197 2419
rect 7019 2312 7053 2346
rect 7091 2312 7125 2346
rect 7163 2312 7197 2346
rect 7019 2239 7053 2273
rect 7091 2239 7125 2273
rect 7163 2239 7197 2273
rect 7019 2166 7053 2200
rect 7091 2166 7125 2200
rect 7163 2166 7197 2200
rect 7019 2092 7053 2126
rect 7091 2092 7125 2126
rect 7163 2092 7197 2126
rect 7019 2018 7053 2052
rect 7091 2018 7125 2052
rect 7163 2018 7197 2052
rect 7019 1944 7053 1978
rect 7091 1944 7125 1978
rect 7163 1944 7197 1978
rect 7019 1870 7053 1904
rect 7091 1870 7125 1904
rect 7163 1870 7197 1904
rect 7019 1796 7053 1830
rect 7091 1796 7125 1830
rect 7163 1796 7197 1830
rect 7019 1722 7053 1756
rect 7091 1722 7125 1756
rect 7163 1722 7197 1756
rect 7019 1648 7053 1682
rect 7091 1648 7125 1682
rect 7163 1648 7197 1682
rect 7019 1574 7053 1608
rect 7091 1574 7125 1608
rect 7163 1574 7197 1608
rect 6840 1144 6946 1250
rect 7587 4092 7621 4118
rect 7515 4082 7693 4092
rect 7515 4048 7519 4082
rect 7519 4048 7587 4082
rect 7587 4048 7621 4082
rect 7621 4048 7689 4082
rect 7689 4048 7693 4082
rect 7515 4014 7693 4048
rect 7515 3980 7519 4014
rect 7519 3980 7587 4014
rect 7587 3980 7621 4014
rect 7621 3980 7689 4014
rect 7689 3980 7693 4014
rect 7515 3946 7693 3980
rect 7515 3912 7519 3946
rect 7519 3912 7587 3946
rect 7587 3912 7621 3946
rect 7621 3912 7689 3946
rect 7689 3912 7693 3946
rect 7515 3878 7693 3912
rect 7515 3844 7519 3878
rect 7519 3844 7587 3878
rect 7587 3844 7621 3878
rect 7621 3844 7689 3878
rect 7689 3844 7693 3878
rect 7515 3810 7693 3844
rect 7515 3776 7519 3810
rect 7519 3776 7587 3810
rect 7587 3776 7621 3810
rect 7621 3776 7689 3810
rect 7689 3776 7693 3810
rect 7515 3742 7693 3776
rect 7515 3708 7519 3742
rect 7519 3708 7587 3742
rect 7587 3708 7621 3742
rect 7621 3708 7689 3742
rect 7689 3708 7693 3742
rect 7515 3674 7693 3708
rect 7515 3640 7519 3674
rect 7519 3640 7587 3674
rect 7587 3640 7621 3674
rect 7621 3640 7689 3674
rect 7689 3640 7693 3674
rect 7515 3606 7693 3640
rect 7515 3572 7519 3606
rect 7519 3572 7587 3606
rect 7587 3572 7621 3606
rect 7621 3572 7689 3606
rect 7689 3572 7693 3606
rect 7515 3538 7693 3572
rect 7515 3504 7519 3538
rect 7519 3504 7587 3538
rect 7587 3504 7621 3538
rect 7621 3504 7689 3538
rect 7689 3504 7693 3538
rect 7515 3470 7693 3504
rect 7515 3436 7519 3470
rect 7519 3436 7587 3470
rect 7587 3436 7621 3470
rect 7621 3436 7689 3470
rect 7689 3436 7693 3470
rect 7515 3402 7693 3436
rect 7515 3368 7519 3402
rect 7519 3368 7587 3402
rect 7587 3368 7621 3402
rect 7621 3368 7689 3402
rect 7689 3368 7693 3402
rect 7515 3334 7693 3368
rect 7515 3300 7519 3334
rect 7519 3300 7587 3334
rect 7587 3300 7621 3334
rect 7621 3300 7689 3334
rect 7689 3300 7693 3334
rect 7515 3266 7693 3300
rect 7515 3232 7519 3266
rect 7519 3232 7587 3266
rect 7587 3232 7621 3266
rect 7621 3232 7689 3266
rect 7689 3232 7693 3266
rect 7515 3198 7693 3232
rect 7515 3194 7519 3198
rect 7519 3194 7587 3198
rect 7587 3194 7621 3198
rect 7621 3194 7689 3198
rect 7689 3194 7693 3198
rect 7587 3164 7621 3182
rect 7587 3148 7621 3164
rect 7515 3074 7549 3108
rect 7587 3074 7621 3108
rect 7659 3074 7693 3108
rect 7515 2994 7549 3028
rect 7587 2994 7621 3028
rect 7659 2994 7693 3028
rect 7515 2914 7549 2948
rect 7587 2914 7621 2948
rect 7659 2914 7693 2948
rect 7515 2834 7549 2868
rect 7587 2834 7621 2868
rect 7659 2834 7693 2868
rect 7515 2754 7549 2788
rect 7587 2754 7621 2788
rect 7659 2754 7693 2788
rect 7515 2674 7549 2708
rect 7587 2674 7621 2708
rect 7659 2674 7693 2708
rect 7515 2594 7549 2628
rect 7587 2594 7621 2628
rect 7659 2594 7693 2628
rect 7587 2540 7621 2556
rect 7587 2522 7621 2540
rect 7515 2506 7519 2518
rect 7519 2506 7587 2518
rect 7587 2506 7621 2518
rect 7621 2506 7689 2518
rect 7689 2506 7693 2518
rect 7515 2472 7693 2506
rect 7515 2438 7519 2472
rect 7519 2438 7587 2472
rect 7587 2438 7621 2472
rect 7621 2438 7689 2472
rect 7689 2438 7693 2472
rect 7515 2404 7693 2438
rect 7515 2370 7519 2404
rect 7519 2370 7587 2404
rect 7587 2370 7621 2404
rect 7621 2370 7689 2404
rect 7689 2370 7693 2404
rect 7515 2336 7693 2370
rect 7515 2302 7519 2336
rect 7519 2302 7587 2336
rect 7587 2302 7621 2336
rect 7621 2302 7689 2336
rect 7689 2302 7693 2336
rect 7515 2268 7693 2302
rect 7515 2234 7519 2268
rect 7519 2234 7587 2268
rect 7587 2234 7621 2268
rect 7621 2234 7689 2268
rect 7689 2234 7693 2268
rect 7515 2200 7693 2234
rect 7515 2166 7519 2200
rect 7519 2166 7587 2200
rect 7587 2166 7621 2200
rect 7621 2166 7689 2200
rect 7689 2166 7693 2200
rect 7515 2132 7693 2166
rect 7515 2098 7519 2132
rect 7519 2098 7587 2132
rect 7587 2098 7621 2132
rect 7621 2098 7689 2132
rect 7689 2098 7693 2132
rect 7515 2064 7693 2098
rect 7515 2030 7519 2064
rect 7519 2030 7587 2064
rect 7587 2030 7621 2064
rect 7621 2030 7689 2064
rect 7689 2030 7693 2064
rect 7515 1996 7693 2030
rect 7515 1962 7519 1996
rect 7519 1962 7587 1996
rect 7587 1962 7621 1996
rect 7621 1962 7689 1996
rect 7689 1962 7693 1996
rect 7515 1928 7693 1962
rect 7515 1894 7519 1928
rect 7519 1894 7587 1928
rect 7587 1894 7621 1928
rect 7621 1894 7689 1928
rect 7689 1894 7693 1928
rect 7515 1860 7693 1894
rect 7515 1826 7519 1860
rect 7519 1826 7587 1860
rect 7587 1826 7621 1860
rect 7621 1826 7689 1860
rect 7689 1826 7693 1860
rect 7515 1792 7693 1826
rect 7515 1758 7519 1792
rect 7519 1758 7587 1792
rect 7587 1758 7621 1792
rect 7621 1758 7689 1792
rect 7689 1758 7693 1792
rect 7515 1724 7693 1758
rect 7515 1690 7519 1724
rect 7519 1690 7587 1724
rect 7587 1690 7621 1724
rect 7621 1690 7689 1724
rect 7689 1690 7693 1724
rect 7515 1656 7693 1690
rect 7515 1622 7519 1656
rect 7519 1622 7587 1656
rect 7587 1622 7621 1656
rect 7621 1622 7689 1656
rect 7689 1622 7693 1656
rect 7515 1620 7693 1622
rect 7587 1586 7621 1620
rect 7270 1144 7376 1250
rect 8011 4064 8045 4098
rect 8083 4064 8117 4098
rect 8155 4064 8189 4098
rect 8011 3991 8045 4025
rect 8083 3991 8117 4025
rect 8155 3991 8189 4025
rect 8011 3918 8045 3952
rect 8083 3918 8117 3952
rect 8155 3918 8189 3952
rect 8011 3845 8045 3879
rect 8083 3845 8117 3879
rect 8155 3845 8189 3879
rect 8011 3772 8045 3806
rect 8083 3772 8117 3806
rect 8155 3772 8189 3806
rect 8011 3699 8045 3733
rect 8083 3699 8117 3733
rect 8155 3699 8189 3733
rect 8011 3626 8045 3660
rect 8083 3626 8117 3660
rect 8155 3626 8189 3660
rect 8011 3553 8045 3587
rect 8083 3553 8117 3587
rect 8155 3553 8189 3587
rect 8011 3480 8045 3514
rect 8083 3480 8117 3514
rect 8155 3480 8189 3514
rect 8011 3407 8045 3441
rect 8083 3407 8117 3441
rect 8155 3407 8189 3441
rect 8011 3334 8045 3368
rect 8083 3334 8117 3368
rect 8155 3334 8189 3368
rect 8011 3261 8045 3295
rect 8083 3261 8117 3295
rect 8155 3261 8189 3295
rect 8011 3188 8045 3222
rect 8083 3188 8117 3222
rect 8155 3188 8189 3222
rect 8011 3115 8045 3149
rect 8083 3115 8117 3149
rect 8155 3115 8189 3149
rect 8011 3042 8045 3076
rect 8083 3042 8117 3076
rect 8155 3042 8189 3076
rect 8011 2969 8045 3003
rect 8083 2969 8117 3003
rect 8155 2969 8189 3003
rect 8011 2896 8045 2930
rect 8083 2896 8117 2930
rect 8155 2896 8189 2930
rect 8011 2823 8045 2857
rect 8083 2823 8117 2857
rect 8155 2823 8189 2857
rect 8011 2750 8045 2784
rect 8083 2750 8117 2784
rect 8155 2750 8189 2784
rect 8011 2677 8045 2711
rect 8083 2677 8117 2711
rect 8155 2677 8189 2711
rect 8011 2604 8045 2638
rect 8083 2604 8117 2638
rect 8155 2604 8189 2638
rect 8011 2531 8045 2565
rect 8083 2531 8117 2565
rect 8155 2531 8189 2565
rect 8011 2458 8045 2492
rect 8083 2458 8117 2492
rect 8155 2458 8189 2492
rect 8011 2385 8045 2419
rect 8083 2385 8117 2419
rect 8155 2385 8189 2419
rect 8011 2312 8045 2346
rect 8083 2312 8117 2346
rect 8155 2312 8189 2346
rect 8011 2239 8045 2273
rect 8083 2239 8117 2273
rect 8155 2239 8189 2273
rect 8011 2166 8045 2200
rect 8083 2166 8117 2200
rect 8155 2166 8189 2200
rect 8011 2092 8045 2126
rect 8083 2092 8117 2126
rect 8155 2092 8189 2126
rect 8011 2018 8045 2052
rect 8083 2018 8117 2052
rect 8155 2018 8189 2052
rect 8011 1944 8045 1978
rect 8083 1944 8117 1978
rect 8155 1944 8189 1978
rect 8011 1870 8045 1904
rect 8083 1870 8117 1904
rect 8155 1870 8189 1904
rect 8011 1796 8045 1830
rect 8083 1796 8117 1830
rect 8155 1796 8189 1830
rect 8011 1722 8045 1756
rect 8083 1722 8117 1756
rect 8155 1722 8189 1756
rect 8011 1648 8045 1682
rect 8083 1648 8117 1682
rect 8155 1648 8189 1682
rect 8011 1574 8045 1608
rect 8083 1574 8117 1608
rect 8155 1574 8189 1608
rect 7832 1144 7938 1250
rect 8579 4092 8613 4118
rect 8507 4082 8685 4092
rect 8507 4048 8511 4082
rect 8511 4048 8579 4082
rect 8579 4048 8613 4082
rect 8613 4048 8681 4082
rect 8681 4048 8685 4082
rect 8507 4014 8685 4048
rect 8507 3980 8511 4014
rect 8511 3980 8579 4014
rect 8579 3980 8613 4014
rect 8613 3980 8681 4014
rect 8681 3980 8685 4014
rect 8507 3946 8685 3980
rect 8507 3912 8511 3946
rect 8511 3912 8579 3946
rect 8579 3912 8613 3946
rect 8613 3912 8681 3946
rect 8681 3912 8685 3946
rect 8507 3878 8685 3912
rect 8507 3844 8511 3878
rect 8511 3844 8579 3878
rect 8579 3844 8613 3878
rect 8613 3844 8681 3878
rect 8681 3844 8685 3878
rect 8507 3810 8685 3844
rect 8507 3776 8511 3810
rect 8511 3776 8579 3810
rect 8579 3776 8613 3810
rect 8613 3776 8681 3810
rect 8681 3776 8685 3810
rect 8507 3742 8685 3776
rect 8507 3708 8511 3742
rect 8511 3708 8579 3742
rect 8579 3708 8613 3742
rect 8613 3708 8681 3742
rect 8681 3708 8685 3742
rect 8507 3674 8685 3708
rect 8507 3640 8511 3674
rect 8511 3640 8579 3674
rect 8579 3640 8613 3674
rect 8613 3640 8681 3674
rect 8681 3640 8685 3674
rect 8507 3606 8685 3640
rect 8507 3572 8511 3606
rect 8511 3572 8579 3606
rect 8579 3572 8613 3606
rect 8613 3572 8681 3606
rect 8681 3572 8685 3606
rect 8507 3538 8685 3572
rect 8507 3504 8511 3538
rect 8511 3504 8579 3538
rect 8579 3504 8613 3538
rect 8613 3504 8681 3538
rect 8681 3504 8685 3538
rect 8507 3470 8685 3504
rect 8507 3436 8511 3470
rect 8511 3436 8579 3470
rect 8579 3436 8613 3470
rect 8613 3436 8681 3470
rect 8681 3436 8685 3470
rect 8507 3402 8685 3436
rect 8507 3368 8511 3402
rect 8511 3368 8579 3402
rect 8579 3368 8613 3402
rect 8613 3368 8681 3402
rect 8681 3368 8685 3402
rect 8507 3334 8685 3368
rect 8507 3300 8511 3334
rect 8511 3300 8579 3334
rect 8579 3300 8613 3334
rect 8613 3300 8681 3334
rect 8681 3300 8685 3334
rect 8507 3266 8685 3300
rect 8507 3232 8511 3266
rect 8511 3232 8579 3266
rect 8579 3232 8613 3266
rect 8613 3232 8681 3266
rect 8681 3232 8685 3266
rect 8507 3198 8685 3232
rect 8507 3194 8511 3198
rect 8511 3194 8579 3198
rect 8579 3194 8613 3198
rect 8613 3194 8681 3198
rect 8681 3194 8685 3198
rect 8579 3164 8613 3182
rect 8579 3148 8613 3164
rect 8507 3074 8541 3108
rect 8579 3074 8613 3108
rect 8651 3074 8685 3108
rect 8507 2994 8541 3028
rect 8579 2994 8613 3028
rect 8651 2994 8685 3028
rect 8507 2914 8541 2948
rect 8579 2914 8613 2948
rect 8651 2914 8685 2948
rect 8507 2834 8541 2868
rect 8579 2834 8613 2868
rect 8651 2834 8685 2868
rect 8507 2754 8541 2788
rect 8579 2754 8613 2788
rect 8651 2754 8685 2788
rect 8507 2674 8541 2708
rect 8579 2674 8613 2708
rect 8651 2674 8685 2708
rect 8507 2594 8541 2628
rect 8579 2594 8613 2628
rect 8651 2594 8685 2628
rect 8579 2540 8613 2556
rect 8579 2522 8613 2540
rect 8507 2506 8511 2518
rect 8511 2506 8579 2518
rect 8579 2506 8613 2518
rect 8613 2506 8681 2518
rect 8681 2506 8685 2518
rect 8507 2472 8685 2506
rect 8507 2438 8511 2472
rect 8511 2438 8579 2472
rect 8579 2438 8613 2472
rect 8613 2438 8681 2472
rect 8681 2438 8685 2472
rect 8507 2404 8685 2438
rect 8507 2370 8511 2404
rect 8511 2370 8579 2404
rect 8579 2370 8613 2404
rect 8613 2370 8681 2404
rect 8681 2370 8685 2404
rect 8507 2336 8685 2370
rect 8507 2302 8511 2336
rect 8511 2302 8579 2336
rect 8579 2302 8613 2336
rect 8613 2302 8681 2336
rect 8681 2302 8685 2336
rect 8507 2268 8685 2302
rect 8507 2234 8511 2268
rect 8511 2234 8579 2268
rect 8579 2234 8613 2268
rect 8613 2234 8681 2268
rect 8681 2234 8685 2268
rect 8507 2200 8685 2234
rect 8507 2166 8511 2200
rect 8511 2166 8579 2200
rect 8579 2166 8613 2200
rect 8613 2166 8681 2200
rect 8681 2166 8685 2200
rect 8507 2132 8685 2166
rect 8507 2098 8511 2132
rect 8511 2098 8579 2132
rect 8579 2098 8613 2132
rect 8613 2098 8681 2132
rect 8681 2098 8685 2132
rect 8507 2064 8685 2098
rect 8507 2030 8511 2064
rect 8511 2030 8579 2064
rect 8579 2030 8613 2064
rect 8613 2030 8681 2064
rect 8681 2030 8685 2064
rect 8507 1996 8685 2030
rect 8507 1962 8511 1996
rect 8511 1962 8579 1996
rect 8579 1962 8613 1996
rect 8613 1962 8681 1996
rect 8681 1962 8685 1996
rect 8507 1928 8685 1962
rect 8507 1894 8511 1928
rect 8511 1894 8579 1928
rect 8579 1894 8613 1928
rect 8613 1894 8681 1928
rect 8681 1894 8685 1928
rect 8507 1860 8685 1894
rect 8507 1826 8511 1860
rect 8511 1826 8579 1860
rect 8579 1826 8613 1860
rect 8613 1826 8681 1860
rect 8681 1826 8685 1860
rect 8507 1792 8685 1826
rect 8507 1758 8511 1792
rect 8511 1758 8579 1792
rect 8579 1758 8613 1792
rect 8613 1758 8681 1792
rect 8681 1758 8685 1792
rect 8507 1724 8685 1758
rect 8507 1690 8511 1724
rect 8511 1690 8579 1724
rect 8579 1690 8613 1724
rect 8613 1690 8681 1724
rect 8681 1690 8685 1724
rect 8507 1656 8685 1690
rect 8507 1622 8511 1656
rect 8511 1622 8579 1656
rect 8579 1622 8613 1656
rect 8613 1622 8681 1656
rect 8681 1622 8685 1656
rect 8507 1620 8685 1622
rect 8579 1586 8613 1620
rect 8262 1144 8368 1250
rect 9003 4064 9037 4098
rect 9075 4064 9109 4098
rect 9147 4064 9181 4098
rect 9003 3991 9037 4025
rect 9075 3991 9109 4025
rect 9147 3991 9181 4025
rect 9003 3918 9037 3952
rect 9075 3918 9109 3952
rect 9147 3918 9181 3952
rect 9003 3845 9037 3879
rect 9075 3845 9109 3879
rect 9147 3845 9181 3879
rect 9003 3772 9037 3806
rect 9075 3772 9109 3806
rect 9147 3772 9181 3806
rect 9003 3699 9037 3733
rect 9075 3699 9109 3733
rect 9147 3699 9181 3733
rect 9003 3626 9037 3660
rect 9075 3626 9109 3660
rect 9147 3626 9181 3660
rect 9003 3553 9037 3587
rect 9075 3553 9109 3587
rect 9147 3553 9181 3587
rect 9003 3480 9037 3514
rect 9075 3480 9109 3514
rect 9147 3480 9181 3514
rect 9003 3407 9037 3441
rect 9075 3407 9109 3441
rect 9147 3407 9181 3441
rect 9003 3334 9037 3368
rect 9075 3334 9109 3368
rect 9147 3334 9181 3368
rect 9003 3261 9037 3295
rect 9075 3261 9109 3295
rect 9147 3261 9181 3295
rect 9003 3188 9037 3222
rect 9075 3188 9109 3222
rect 9147 3188 9181 3222
rect 9003 3115 9037 3149
rect 9075 3115 9109 3149
rect 9147 3115 9181 3149
rect 9003 3042 9037 3076
rect 9075 3042 9109 3076
rect 9147 3042 9181 3076
rect 9003 2969 9037 3003
rect 9075 2969 9109 3003
rect 9147 2969 9181 3003
rect 9003 2896 9037 2930
rect 9075 2896 9109 2930
rect 9147 2896 9181 2930
rect 9003 2823 9037 2857
rect 9075 2823 9109 2857
rect 9147 2823 9181 2857
rect 9003 2750 9037 2784
rect 9075 2750 9109 2784
rect 9147 2750 9181 2784
rect 9003 2677 9037 2711
rect 9075 2677 9109 2711
rect 9147 2677 9181 2711
rect 9003 2604 9037 2638
rect 9075 2604 9109 2638
rect 9147 2604 9181 2638
rect 9003 2531 9037 2565
rect 9075 2531 9109 2565
rect 9147 2531 9181 2565
rect 9003 2458 9037 2492
rect 9075 2458 9109 2492
rect 9147 2458 9181 2492
rect 9003 2385 9037 2419
rect 9075 2385 9109 2419
rect 9147 2385 9181 2419
rect 9003 2312 9037 2346
rect 9075 2312 9109 2346
rect 9147 2312 9181 2346
rect 9003 2239 9037 2273
rect 9075 2239 9109 2273
rect 9147 2239 9181 2273
rect 9003 2166 9037 2200
rect 9075 2166 9109 2200
rect 9147 2166 9181 2200
rect 9003 2092 9037 2126
rect 9075 2092 9109 2126
rect 9147 2092 9181 2126
rect 9003 2018 9037 2052
rect 9075 2018 9109 2052
rect 9147 2018 9181 2052
rect 9003 1944 9037 1978
rect 9075 1944 9109 1978
rect 9147 1944 9181 1978
rect 9003 1870 9037 1904
rect 9075 1870 9109 1904
rect 9147 1870 9181 1904
rect 9003 1796 9037 1830
rect 9075 1796 9109 1830
rect 9147 1796 9181 1830
rect 9003 1722 9037 1756
rect 9075 1722 9109 1756
rect 9147 1722 9181 1756
rect 9003 1648 9037 1682
rect 9075 1648 9109 1682
rect 9147 1648 9181 1682
rect 9003 1574 9037 1608
rect 9075 1574 9109 1608
rect 9147 1574 9181 1608
rect 8824 1144 8930 1250
rect 9571 4092 9605 4118
rect 9499 4082 9677 4092
rect 9499 4048 9503 4082
rect 9503 4048 9571 4082
rect 9571 4048 9605 4082
rect 9605 4048 9673 4082
rect 9673 4048 9677 4082
rect 9499 4014 9677 4048
rect 9499 3980 9503 4014
rect 9503 3980 9571 4014
rect 9571 3980 9605 4014
rect 9605 3980 9673 4014
rect 9673 3980 9677 4014
rect 9499 3946 9677 3980
rect 9499 3912 9503 3946
rect 9503 3912 9571 3946
rect 9571 3912 9605 3946
rect 9605 3912 9673 3946
rect 9673 3912 9677 3946
rect 9499 3878 9677 3912
rect 9499 3844 9503 3878
rect 9503 3844 9571 3878
rect 9571 3844 9605 3878
rect 9605 3844 9673 3878
rect 9673 3844 9677 3878
rect 9499 3810 9677 3844
rect 9499 3776 9503 3810
rect 9503 3776 9571 3810
rect 9571 3776 9605 3810
rect 9605 3776 9673 3810
rect 9673 3776 9677 3810
rect 9499 3742 9677 3776
rect 9499 3708 9503 3742
rect 9503 3708 9571 3742
rect 9571 3708 9605 3742
rect 9605 3708 9673 3742
rect 9673 3708 9677 3742
rect 9499 3674 9677 3708
rect 9499 3640 9503 3674
rect 9503 3640 9571 3674
rect 9571 3640 9605 3674
rect 9605 3640 9673 3674
rect 9673 3640 9677 3674
rect 9499 3606 9677 3640
rect 9499 3572 9503 3606
rect 9503 3572 9571 3606
rect 9571 3572 9605 3606
rect 9605 3572 9673 3606
rect 9673 3572 9677 3606
rect 9499 3538 9677 3572
rect 9499 3504 9503 3538
rect 9503 3504 9571 3538
rect 9571 3504 9605 3538
rect 9605 3504 9673 3538
rect 9673 3504 9677 3538
rect 9499 3470 9677 3504
rect 9499 3436 9503 3470
rect 9503 3436 9571 3470
rect 9571 3436 9605 3470
rect 9605 3436 9673 3470
rect 9673 3436 9677 3470
rect 9499 3402 9677 3436
rect 9499 3368 9503 3402
rect 9503 3368 9571 3402
rect 9571 3368 9605 3402
rect 9605 3368 9673 3402
rect 9673 3368 9677 3402
rect 9499 3334 9677 3368
rect 9499 3300 9503 3334
rect 9503 3300 9571 3334
rect 9571 3300 9605 3334
rect 9605 3300 9673 3334
rect 9673 3300 9677 3334
rect 9499 3266 9677 3300
rect 9499 3232 9503 3266
rect 9503 3232 9571 3266
rect 9571 3232 9605 3266
rect 9605 3232 9673 3266
rect 9673 3232 9677 3266
rect 9499 3198 9677 3232
rect 9499 3194 9503 3198
rect 9503 3194 9571 3198
rect 9571 3194 9605 3198
rect 9605 3194 9673 3198
rect 9673 3194 9677 3198
rect 9571 3164 9605 3182
rect 9571 3148 9605 3164
rect 9499 3074 9533 3108
rect 9571 3074 9605 3108
rect 9643 3074 9677 3108
rect 9499 2994 9533 3028
rect 9571 2994 9605 3028
rect 9643 2994 9677 3028
rect 9499 2914 9533 2948
rect 9571 2914 9605 2948
rect 9643 2914 9677 2948
rect 9499 2834 9533 2868
rect 9571 2834 9605 2868
rect 9643 2834 9677 2868
rect 9499 2754 9533 2788
rect 9571 2754 9605 2788
rect 9643 2754 9677 2788
rect 9499 2674 9533 2708
rect 9571 2674 9605 2708
rect 9643 2674 9677 2708
rect 9499 2594 9533 2628
rect 9571 2594 9605 2628
rect 9643 2594 9677 2628
rect 9571 2540 9605 2556
rect 9571 2522 9605 2540
rect 9499 2506 9503 2518
rect 9503 2506 9571 2518
rect 9571 2506 9605 2518
rect 9605 2506 9673 2518
rect 9673 2506 9677 2518
rect 9499 2472 9677 2506
rect 9499 2438 9503 2472
rect 9503 2438 9571 2472
rect 9571 2438 9605 2472
rect 9605 2438 9673 2472
rect 9673 2438 9677 2472
rect 9499 2404 9677 2438
rect 9499 2370 9503 2404
rect 9503 2370 9571 2404
rect 9571 2370 9605 2404
rect 9605 2370 9673 2404
rect 9673 2370 9677 2404
rect 9499 2336 9677 2370
rect 9499 2302 9503 2336
rect 9503 2302 9571 2336
rect 9571 2302 9605 2336
rect 9605 2302 9673 2336
rect 9673 2302 9677 2336
rect 9499 2268 9677 2302
rect 9499 2234 9503 2268
rect 9503 2234 9571 2268
rect 9571 2234 9605 2268
rect 9605 2234 9673 2268
rect 9673 2234 9677 2268
rect 9499 2200 9677 2234
rect 9499 2166 9503 2200
rect 9503 2166 9571 2200
rect 9571 2166 9605 2200
rect 9605 2166 9673 2200
rect 9673 2166 9677 2200
rect 9499 2132 9677 2166
rect 9499 2098 9503 2132
rect 9503 2098 9571 2132
rect 9571 2098 9605 2132
rect 9605 2098 9673 2132
rect 9673 2098 9677 2132
rect 9499 2064 9677 2098
rect 9499 2030 9503 2064
rect 9503 2030 9571 2064
rect 9571 2030 9605 2064
rect 9605 2030 9673 2064
rect 9673 2030 9677 2064
rect 9499 1996 9677 2030
rect 9499 1962 9503 1996
rect 9503 1962 9571 1996
rect 9571 1962 9605 1996
rect 9605 1962 9673 1996
rect 9673 1962 9677 1996
rect 9499 1928 9677 1962
rect 9499 1894 9503 1928
rect 9503 1894 9571 1928
rect 9571 1894 9605 1928
rect 9605 1894 9673 1928
rect 9673 1894 9677 1928
rect 9499 1860 9677 1894
rect 9499 1826 9503 1860
rect 9503 1826 9571 1860
rect 9571 1826 9605 1860
rect 9605 1826 9673 1860
rect 9673 1826 9677 1860
rect 9499 1792 9677 1826
rect 9499 1758 9503 1792
rect 9503 1758 9571 1792
rect 9571 1758 9605 1792
rect 9605 1758 9673 1792
rect 9673 1758 9677 1792
rect 9499 1724 9677 1758
rect 9499 1690 9503 1724
rect 9503 1690 9571 1724
rect 9571 1690 9605 1724
rect 9605 1690 9673 1724
rect 9673 1690 9677 1724
rect 9499 1656 9677 1690
rect 9499 1622 9503 1656
rect 9503 1622 9571 1656
rect 9571 1622 9605 1656
rect 9605 1622 9673 1656
rect 9673 1622 9677 1656
rect 9499 1620 9677 1622
rect 9571 1586 9605 1620
rect 9254 1144 9360 1250
rect 9995 4064 10029 4098
rect 10067 4064 10101 4098
rect 10139 4064 10173 4098
rect 9995 3991 10029 4025
rect 10067 3991 10101 4025
rect 10139 3991 10173 4025
rect 9995 3918 10029 3952
rect 10067 3918 10101 3952
rect 10139 3918 10173 3952
rect 9995 3845 10029 3879
rect 10067 3845 10101 3879
rect 10139 3845 10173 3879
rect 9995 3772 10029 3806
rect 10067 3772 10101 3806
rect 10139 3772 10173 3806
rect 9995 3699 10029 3733
rect 10067 3699 10101 3733
rect 10139 3699 10173 3733
rect 9995 3626 10029 3660
rect 10067 3626 10101 3660
rect 10139 3626 10173 3660
rect 9995 3553 10029 3587
rect 10067 3553 10101 3587
rect 10139 3553 10173 3587
rect 9995 3480 10029 3514
rect 10067 3480 10101 3514
rect 10139 3480 10173 3514
rect 9995 3407 10029 3441
rect 10067 3407 10101 3441
rect 10139 3407 10173 3441
rect 9995 3334 10029 3368
rect 10067 3334 10101 3368
rect 10139 3334 10173 3368
rect 9995 3261 10029 3295
rect 10067 3261 10101 3295
rect 10139 3261 10173 3295
rect 9995 3188 10029 3222
rect 10067 3188 10101 3222
rect 10139 3188 10173 3222
rect 9995 3115 10029 3149
rect 10067 3115 10101 3149
rect 10139 3115 10173 3149
rect 9995 3042 10029 3076
rect 10067 3042 10101 3076
rect 10139 3042 10173 3076
rect 9995 2969 10029 3003
rect 10067 2969 10101 3003
rect 10139 2969 10173 3003
rect 9995 2896 10029 2930
rect 10067 2896 10101 2930
rect 10139 2896 10173 2930
rect 9995 2823 10029 2857
rect 10067 2823 10101 2857
rect 10139 2823 10173 2857
rect 9995 2750 10029 2784
rect 10067 2750 10101 2784
rect 10139 2750 10173 2784
rect 9995 2677 10029 2711
rect 10067 2677 10101 2711
rect 10139 2677 10173 2711
rect 9995 2604 10029 2638
rect 10067 2604 10101 2638
rect 10139 2604 10173 2638
rect 9995 2531 10029 2565
rect 10067 2531 10101 2565
rect 10139 2531 10173 2565
rect 9995 2458 10029 2492
rect 10067 2458 10101 2492
rect 10139 2458 10173 2492
rect 9995 2385 10029 2419
rect 10067 2385 10101 2419
rect 10139 2385 10173 2419
rect 9995 2312 10029 2346
rect 10067 2312 10101 2346
rect 10139 2312 10173 2346
rect 9995 2239 10029 2273
rect 10067 2239 10101 2273
rect 10139 2239 10173 2273
rect 9995 2166 10029 2200
rect 10067 2166 10101 2200
rect 10139 2166 10173 2200
rect 9995 2092 10029 2126
rect 10067 2092 10101 2126
rect 10139 2092 10173 2126
rect 9995 2018 10029 2052
rect 10067 2018 10101 2052
rect 10139 2018 10173 2052
rect 9995 1944 10029 1978
rect 10067 1944 10101 1978
rect 10139 1944 10173 1978
rect 9995 1870 10029 1904
rect 10067 1870 10101 1904
rect 10139 1870 10173 1904
rect 9995 1796 10029 1830
rect 10067 1796 10101 1830
rect 10139 1796 10173 1830
rect 9995 1722 10029 1756
rect 10067 1722 10101 1756
rect 10139 1722 10173 1756
rect 9995 1648 10029 1682
rect 10067 1648 10101 1682
rect 10139 1648 10173 1682
rect 9995 1574 10029 1608
rect 10067 1574 10101 1608
rect 10139 1574 10173 1608
rect 9816 1144 9922 1250
rect 10563 4092 10597 4118
rect 10491 4082 10669 4092
rect 10491 4048 10495 4082
rect 10495 4048 10563 4082
rect 10563 4048 10597 4082
rect 10597 4048 10665 4082
rect 10665 4048 10669 4082
rect 10491 4014 10669 4048
rect 10491 3980 10495 4014
rect 10495 3980 10563 4014
rect 10563 3980 10597 4014
rect 10597 3980 10665 4014
rect 10665 3980 10669 4014
rect 10491 3946 10669 3980
rect 10491 3912 10495 3946
rect 10495 3912 10563 3946
rect 10563 3912 10597 3946
rect 10597 3912 10665 3946
rect 10665 3912 10669 3946
rect 10491 3878 10669 3912
rect 10491 3844 10495 3878
rect 10495 3844 10563 3878
rect 10563 3844 10597 3878
rect 10597 3844 10665 3878
rect 10665 3844 10669 3878
rect 10491 3810 10669 3844
rect 10491 3776 10495 3810
rect 10495 3776 10563 3810
rect 10563 3776 10597 3810
rect 10597 3776 10665 3810
rect 10665 3776 10669 3810
rect 10491 3742 10669 3776
rect 10491 3708 10495 3742
rect 10495 3708 10563 3742
rect 10563 3708 10597 3742
rect 10597 3708 10665 3742
rect 10665 3708 10669 3742
rect 10491 3674 10669 3708
rect 10491 3640 10495 3674
rect 10495 3640 10563 3674
rect 10563 3640 10597 3674
rect 10597 3640 10665 3674
rect 10665 3640 10669 3674
rect 10491 3606 10669 3640
rect 10491 3572 10495 3606
rect 10495 3572 10563 3606
rect 10563 3572 10597 3606
rect 10597 3572 10665 3606
rect 10665 3572 10669 3606
rect 10491 3538 10669 3572
rect 10491 3504 10495 3538
rect 10495 3504 10563 3538
rect 10563 3504 10597 3538
rect 10597 3504 10665 3538
rect 10665 3504 10669 3538
rect 10491 3470 10669 3504
rect 10491 3436 10495 3470
rect 10495 3436 10563 3470
rect 10563 3436 10597 3470
rect 10597 3436 10665 3470
rect 10665 3436 10669 3470
rect 10491 3402 10669 3436
rect 10491 3368 10495 3402
rect 10495 3368 10563 3402
rect 10563 3368 10597 3402
rect 10597 3368 10665 3402
rect 10665 3368 10669 3402
rect 10491 3334 10669 3368
rect 10491 3300 10495 3334
rect 10495 3300 10563 3334
rect 10563 3300 10597 3334
rect 10597 3300 10665 3334
rect 10665 3300 10669 3334
rect 10491 3266 10669 3300
rect 10491 3232 10495 3266
rect 10495 3232 10563 3266
rect 10563 3232 10597 3266
rect 10597 3232 10665 3266
rect 10665 3232 10669 3266
rect 10491 3198 10669 3232
rect 10491 3194 10495 3198
rect 10495 3194 10563 3198
rect 10563 3194 10597 3198
rect 10597 3194 10665 3198
rect 10665 3194 10669 3198
rect 10563 3164 10597 3182
rect 10563 3148 10597 3164
rect 10491 3074 10525 3108
rect 10563 3074 10597 3108
rect 10635 3074 10669 3108
rect 10491 2994 10525 3028
rect 10563 2994 10597 3028
rect 10635 2994 10669 3028
rect 10491 2914 10525 2948
rect 10563 2914 10597 2948
rect 10635 2914 10669 2948
rect 10491 2834 10525 2868
rect 10563 2834 10597 2868
rect 10635 2834 10669 2868
rect 10491 2754 10525 2788
rect 10563 2754 10597 2788
rect 10635 2754 10669 2788
rect 10491 2674 10525 2708
rect 10563 2674 10597 2708
rect 10635 2674 10669 2708
rect 10491 2594 10525 2628
rect 10563 2594 10597 2628
rect 10635 2594 10669 2628
rect 10563 2540 10597 2556
rect 10563 2522 10597 2540
rect 10491 2506 10495 2518
rect 10495 2506 10563 2518
rect 10563 2506 10597 2518
rect 10597 2506 10665 2518
rect 10665 2506 10669 2518
rect 10491 2472 10669 2506
rect 10491 2438 10495 2472
rect 10495 2438 10563 2472
rect 10563 2438 10597 2472
rect 10597 2438 10665 2472
rect 10665 2438 10669 2472
rect 10491 2404 10669 2438
rect 10491 2370 10495 2404
rect 10495 2370 10563 2404
rect 10563 2370 10597 2404
rect 10597 2370 10665 2404
rect 10665 2370 10669 2404
rect 10491 2336 10669 2370
rect 10491 2302 10495 2336
rect 10495 2302 10563 2336
rect 10563 2302 10597 2336
rect 10597 2302 10665 2336
rect 10665 2302 10669 2336
rect 10491 2268 10669 2302
rect 10491 2234 10495 2268
rect 10495 2234 10563 2268
rect 10563 2234 10597 2268
rect 10597 2234 10665 2268
rect 10665 2234 10669 2268
rect 10491 2200 10669 2234
rect 10491 2166 10495 2200
rect 10495 2166 10563 2200
rect 10563 2166 10597 2200
rect 10597 2166 10665 2200
rect 10665 2166 10669 2200
rect 10491 2132 10669 2166
rect 10491 2098 10495 2132
rect 10495 2098 10563 2132
rect 10563 2098 10597 2132
rect 10597 2098 10665 2132
rect 10665 2098 10669 2132
rect 10491 2064 10669 2098
rect 10491 2030 10495 2064
rect 10495 2030 10563 2064
rect 10563 2030 10597 2064
rect 10597 2030 10665 2064
rect 10665 2030 10669 2064
rect 10491 1996 10669 2030
rect 10491 1962 10495 1996
rect 10495 1962 10563 1996
rect 10563 1962 10597 1996
rect 10597 1962 10665 1996
rect 10665 1962 10669 1996
rect 10491 1928 10669 1962
rect 10491 1894 10495 1928
rect 10495 1894 10563 1928
rect 10563 1894 10597 1928
rect 10597 1894 10665 1928
rect 10665 1894 10669 1928
rect 10491 1860 10669 1894
rect 10491 1826 10495 1860
rect 10495 1826 10563 1860
rect 10563 1826 10597 1860
rect 10597 1826 10665 1860
rect 10665 1826 10669 1860
rect 10491 1792 10669 1826
rect 10491 1758 10495 1792
rect 10495 1758 10563 1792
rect 10563 1758 10597 1792
rect 10597 1758 10665 1792
rect 10665 1758 10669 1792
rect 10491 1724 10669 1758
rect 10491 1690 10495 1724
rect 10495 1690 10563 1724
rect 10563 1690 10597 1724
rect 10597 1690 10665 1724
rect 10665 1690 10669 1724
rect 10491 1656 10669 1690
rect 10491 1622 10495 1656
rect 10495 1622 10563 1656
rect 10563 1622 10597 1656
rect 10597 1622 10665 1656
rect 10665 1622 10669 1656
rect 10491 1620 10669 1622
rect 10563 1586 10597 1620
rect 10246 1144 10352 1250
rect 10987 4064 11021 4098
rect 11059 4064 11093 4098
rect 11131 4064 11165 4098
rect 10987 3991 11021 4025
rect 11059 3991 11093 4025
rect 11131 3991 11165 4025
rect 10987 3918 11021 3952
rect 11059 3918 11093 3952
rect 11131 3918 11165 3952
rect 10987 3845 11021 3879
rect 11059 3845 11093 3879
rect 11131 3845 11165 3879
rect 10987 3772 11021 3806
rect 11059 3772 11093 3806
rect 11131 3772 11165 3806
rect 10987 3699 11021 3733
rect 11059 3699 11093 3733
rect 11131 3699 11165 3733
rect 10987 3626 11021 3660
rect 11059 3626 11093 3660
rect 11131 3626 11165 3660
rect 10987 3553 11021 3587
rect 11059 3553 11093 3587
rect 11131 3553 11165 3587
rect 10987 3480 11021 3514
rect 11059 3480 11093 3514
rect 11131 3480 11165 3514
rect 10987 3407 11021 3441
rect 11059 3407 11093 3441
rect 11131 3407 11165 3441
rect 10987 3334 11021 3368
rect 11059 3334 11093 3368
rect 11131 3334 11165 3368
rect 10987 3261 11021 3295
rect 11059 3261 11093 3295
rect 11131 3261 11165 3295
rect 10987 3188 11021 3222
rect 11059 3188 11093 3222
rect 11131 3188 11165 3222
rect 10987 3115 11021 3149
rect 11059 3115 11093 3149
rect 11131 3115 11165 3149
rect 10987 3042 11021 3076
rect 11059 3042 11093 3076
rect 11131 3042 11165 3076
rect 10987 2969 11021 3003
rect 11059 2969 11093 3003
rect 11131 2969 11165 3003
rect 10987 2896 11021 2930
rect 11059 2896 11093 2930
rect 11131 2896 11165 2930
rect 10987 2823 11021 2857
rect 11059 2823 11093 2857
rect 11131 2823 11165 2857
rect 10987 2750 11021 2784
rect 11059 2750 11093 2784
rect 11131 2750 11165 2784
rect 10987 2677 11021 2711
rect 11059 2677 11093 2711
rect 11131 2677 11165 2711
rect 10987 2604 11021 2638
rect 11059 2604 11093 2638
rect 11131 2604 11165 2638
rect 10987 2531 11021 2565
rect 11059 2531 11093 2565
rect 11131 2531 11165 2565
rect 10987 2458 11021 2492
rect 11059 2458 11093 2492
rect 11131 2458 11165 2492
rect 10987 2385 11021 2419
rect 11059 2385 11093 2419
rect 11131 2385 11165 2419
rect 10987 2312 11021 2346
rect 11059 2312 11093 2346
rect 11131 2312 11165 2346
rect 10987 2239 11021 2273
rect 11059 2239 11093 2273
rect 11131 2239 11165 2273
rect 10987 2166 11021 2200
rect 11059 2166 11093 2200
rect 11131 2166 11165 2200
rect 10987 2092 11021 2126
rect 11059 2092 11093 2126
rect 11131 2092 11165 2126
rect 10987 2018 11021 2052
rect 11059 2018 11093 2052
rect 11131 2018 11165 2052
rect 10987 1944 11021 1978
rect 11059 1944 11093 1978
rect 11131 1944 11165 1978
rect 10987 1870 11021 1904
rect 11059 1870 11093 1904
rect 11131 1870 11165 1904
rect 10987 1796 11021 1830
rect 11059 1796 11093 1830
rect 11131 1796 11165 1830
rect 10987 1722 11021 1756
rect 11059 1722 11093 1756
rect 11131 1722 11165 1756
rect 10987 1648 11021 1682
rect 11059 1648 11093 1682
rect 11131 1648 11165 1682
rect 10987 1574 11021 1608
rect 11059 1574 11093 1608
rect 11131 1574 11165 1608
rect 10808 1144 10914 1250
rect 11555 4092 11589 4118
rect 11483 4082 11661 4092
rect 11483 4048 11487 4082
rect 11487 4048 11555 4082
rect 11555 4048 11589 4082
rect 11589 4048 11657 4082
rect 11657 4048 11661 4082
rect 11483 4014 11661 4048
rect 11483 3980 11487 4014
rect 11487 3980 11555 4014
rect 11555 3980 11589 4014
rect 11589 3980 11657 4014
rect 11657 3980 11661 4014
rect 11483 3946 11661 3980
rect 11483 3912 11487 3946
rect 11487 3912 11555 3946
rect 11555 3912 11589 3946
rect 11589 3912 11657 3946
rect 11657 3912 11661 3946
rect 11483 3878 11661 3912
rect 11483 3844 11487 3878
rect 11487 3844 11555 3878
rect 11555 3844 11589 3878
rect 11589 3844 11657 3878
rect 11657 3844 11661 3878
rect 11483 3810 11661 3844
rect 11483 3776 11487 3810
rect 11487 3776 11555 3810
rect 11555 3776 11589 3810
rect 11589 3776 11657 3810
rect 11657 3776 11661 3810
rect 11483 3742 11661 3776
rect 11483 3708 11487 3742
rect 11487 3708 11555 3742
rect 11555 3708 11589 3742
rect 11589 3708 11657 3742
rect 11657 3708 11661 3742
rect 11483 3674 11661 3708
rect 11483 3640 11487 3674
rect 11487 3640 11555 3674
rect 11555 3640 11589 3674
rect 11589 3640 11657 3674
rect 11657 3640 11661 3674
rect 11483 3606 11661 3640
rect 11483 3572 11487 3606
rect 11487 3572 11555 3606
rect 11555 3572 11589 3606
rect 11589 3572 11657 3606
rect 11657 3572 11661 3606
rect 11483 3538 11661 3572
rect 11483 3504 11487 3538
rect 11487 3504 11555 3538
rect 11555 3504 11589 3538
rect 11589 3504 11657 3538
rect 11657 3504 11661 3538
rect 11483 3470 11661 3504
rect 11483 3436 11487 3470
rect 11487 3436 11555 3470
rect 11555 3436 11589 3470
rect 11589 3436 11657 3470
rect 11657 3436 11661 3470
rect 11483 3402 11661 3436
rect 11483 3368 11487 3402
rect 11487 3368 11555 3402
rect 11555 3368 11589 3402
rect 11589 3368 11657 3402
rect 11657 3368 11661 3402
rect 11483 3334 11661 3368
rect 11483 3300 11487 3334
rect 11487 3300 11555 3334
rect 11555 3300 11589 3334
rect 11589 3300 11657 3334
rect 11657 3300 11661 3334
rect 11483 3266 11661 3300
rect 11483 3232 11487 3266
rect 11487 3232 11555 3266
rect 11555 3232 11589 3266
rect 11589 3232 11657 3266
rect 11657 3232 11661 3266
rect 11483 3198 11661 3232
rect 11483 3194 11487 3198
rect 11487 3194 11555 3198
rect 11555 3194 11589 3198
rect 11589 3194 11657 3198
rect 11657 3194 11661 3198
rect 11555 3164 11589 3182
rect 11555 3148 11589 3164
rect 11483 3074 11517 3108
rect 11555 3074 11589 3108
rect 11627 3074 11661 3108
rect 11483 2994 11517 3028
rect 11555 2994 11589 3028
rect 11627 2994 11661 3028
rect 11483 2914 11517 2948
rect 11555 2914 11589 2948
rect 11627 2914 11661 2948
rect 11483 2834 11517 2868
rect 11555 2834 11589 2868
rect 11627 2834 11661 2868
rect 11483 2754 11517 2788
rect 11555 2754 11589 2788
rect 11627 2754 11661 2788
rect 11483 2674 11517 2708
rect 11555 2674 11589 2708
rect 11627 2674 11661 2708
rect 11483 2594 11517 2628
rect 11555 2594 11589 2628
rect 11627 2594 11661 2628
rect 11555 2540 11589 2556
rect 11555 2522 11589 2540
rect 11483 2506 11487 2518
rect 11487 2506 11555 2518
rect 11555 2506 11589 2518
rect 11589 2506 11657 2518
rect 11657 2506 11661 2518
rect 11483 2472 11661 2506
rect 11483 2438 11487 2472
rect 11487 2438 11555 2472
rect 11555 2438 11589 2472
rect 11589 2438 11657 2472
rect 11657 2438 11661 2472
rect 11483 2404 11661 2438
rect 11483 2370 11487 2404
rect 11487 2370 11555 2404
rect 11555 2370 11589 2404
rect 11589 2370 11657 2404
rect 11657 2370 11661 2404
rect 11483 2336 11661 2370
rect 11483 2302 11487 2336
rect 11487 2302 11555 2336
rect 11555 2302 11589 2336
rect 11589 2302 11657 2336
rect 11657 2302 11661 2336
rect 11483 2268 11661 2302
rect 11483 2234 11487 2268
rect 11487 2234 11555 2268
rect 11555 2234 11589 2268
rect 11589 2234 11657 2268
rect 11657 2234 11661 2268
rect 11483 2200 11661 2234
rect 11483 2166 11487 2200
rect 11487 2166 11555 2200
rect 11555 2166 11589 2200
rect 11589 2166 11657 2200
rect 11657 2166 11661 2200
rect 11483 2132 11661 2166
rect 11483 2098 11487 2132
rect 11487 2098 11555 2132
rect 11555 2098 11589 2132
rect 11589 2098 11657 2132
rect 11657 2098 11661 2132
rect 11483 2064 11661 2098
rect 11483 2030 11487 2064
rect 11487 2030 11555 2064
rect 11555 2030 11589 2064
rect 11589 2030 11657 2064
rect 11657 2030 11661 2064
rect 11483 1996 11661 2030
rect 11483 1962 11487 1996
rect 11487 1962 11555 1996
rect 11555 1962 11589 1996
rect 11589 1962 11657 1996
rect 11657 1962 11661 1996
rect 11483 1928 11661 1962
rect 11483 1894 11487 1928
rect 11487 1894 11555 1928
rect 11555 1894 11589 1928
rect 11589 1894 11657 1928
rect 11657 1894 11661 1928
rect 11483 1860 11661 1894
rect 11483 1826 11487 1860
rect 11487 1826 11555 1860
rect 11555 1826 11589 1860
rect 11589 1826 11657 1860
rect 11657 1826 11661 1860
rect 11483 1792 11661 1826
rect 11483 1758 11487 1792
rect 11487 1758 11555 1792
rect 11555 1758 11589 1792
rect 11589 1758 11657 1792
rect 11657 1758 11661 1792
rect 11483 1724 11661 1758
rect 11483 1690 11487 1724
rect 11487 1690 11555 1724
rect 11555 1690 11589 1724
rect 11589 1690 11657 1724
rect 11657 1690 11661 1724
rect 11483 1656 11661 1690
rect 11483 1622 11487 1656
rect 11487 1622 11555 1656
rect 11555 1622 11589 1656
rect 11589 1622 11657 1656
rect 11657 1622 11661 1656
rect 11483 1620 11661 1622
rect 11555 1586 11589 1620
rect 11238 1144 11344 1250
rect 11979 4064 12013 4098
rect 12051 4064 12085 4098
rect 12123 4064 12157 4098
rect 11979 3991 12013 4025
rect 12051 3991 12085 4025
rect 12123 3991 12157 4025
rect 11979 3918 12013 3952
rect 12051 3918 12085 3952
rect 12123 3918 12157 3952
rect 11979 3845 12013 3879
rect 12051 3845 12085 3879
rect 12123 3845 12157 3879
rect 11979 3772 12013 3806
rect 12051 3772 12085 3806
rect 12123 3772 12157 3806
rect 11979 3699 12013 3733
rect 12051 3699 12085 3733
rect 12123 3699 12157 3733
rect 11979 3626 12013 3660
rect 12051 3626 12085 3660
rect 12123 3626 12157 3660
rect 11979 3553 12013 3587
rect 12051 3553 12085 3587
rect 12123 3553 12157 3587
rect 11979 3480 12013 3514
rect 12051 3480 12085 3514
rect 12123 3480 12157 3514
rect 11979 3407 12013 3441
rect 12051 3407 12085 3441
rect 12123 3407 12157 3441
rect 11979 3334 12013 3368
rect 12051 3334 12085 3368
rect 12123 3334 12157 3368
rect 11979 3261 12013 3295
rect 12051 3261 12085 3295
rect 12123 3261 12157 3295
rect 11979 3188 12013 3222
rect 12051 3188 12085 3222
rect 12123 3188 12157 3222
rect 11979 3115 12013 3149
rect 12051 3115 12085 3149
rect 12123 3115 12157 3149
rect 11979 3042 12013 3076
rect 12051 3042 12085 3076
rect 12123 3042 12157 3076
rect 11979 2969 12013 3003
rect 12051 2969 12085 3003
rect 12123 2969 12157 3003
rect 11979 2896 12013 2930
rect 12051 2896 12085 2930
rect 12123 2896 12157 2930
rect 11979 2823 12013 2857
rect 12051 2823 12085 2857
rect 12123 2823 12157 2857
rect 11979 2750 12013 2784
rect 12051 2750 12085 2784
rect 12123 2750 12157 2784
rect 11979 2677 12013 2711
rect 12051 2677 12085 2711
rect 12123 2677 12157 2711
rect 11979 2604 12013 2638
rect 12051 2604 12085 2638
rect 12123 2604 12157 2638
rect 11979 2531 12013 2565
rect 12051 2531 12085 2565
rect 12123 2531 12157 2565
rect 11979 2458 12013 2492
rect 12051 2458 12085 2492
rect 12123 2458 12157 2492
rect 11979 2385 12013 2419
rect 12051 2385 12085 2419
rect 12123 2385 12157 2419
rect 11979 2312 12013 2346
rect 12051 2312 12085 2346
rect 12123 2312 12157 2346
rect 11979 2239 12013 2273
rect 12051 2239 12085 2273
rect 12123 2239 12157 2273
rect 11979 2166 12013 2200
rect 12051 2166 12085 2200
rect 12123 2166 12157 2200
rect 11979 2092 12013 2126
rect 12051 2092 12085 2126
rect 12123 2092 12157 2126
rect 11979 2018 12013 2052
rect 12051 2018 12085 2052
rect 12123 2018 12157 2052
rect 11979 1944 12013 1978
rect 12051 1944 12085 1978
rect 12123 1944 12157 1978
rect 11979 1870 12013 1904
rect 12051 1870 12085 1904
rect 12123 1870 12157 1904
rect 11979 1796 12013 1830
rect 12051 1796 12085 1830
rect 12123 1796 12157 1830
rect 11979 1722 12013 1756
rect 12051 1722 12085 1756
rect 12123 1722 12157 1756
rect 11979 1648 12013 1682
rect 12051 1648 12085 1682
rect 12123 1648 12157 1682
rect 11979 1574 12013 1608
rect 12051 1574 12085 1608
rect 12123 1574 12157 1608
rect 11800 1144 11906 1250
rect 12547 4092 12581 4118
rect 12475 4082 12653 4092
rect 12475 4048 12479 4082
rect 12479 4048 12547 4082
rect 12547 4048 12581 4082
rect 12581 4048 12649 4082
rect 12649 4048 12653 4082
rect 12475 4014 12653 4048
rect 12475 3980 12479 4014
rect 12479 3980 12547 4014
rect 12547 3980 12581 4014
rect 12581 3980 12649 4014
rect 12649 3980 12653 4014
rect 12475 3946 12653 3980
rect 12475 3912 12479 3946
rect 12479 3912 12547 3946
rect 12547 3912 12581 3946
rect 12581 3912 12649 3946
rect 12649 3912 12653 3946
rect 12475 3878 12653 3912
rect 12475 3844 12479 3878
rect 12479 3844 12547 3878
rect 12547 3844 12581 3878
rect 12581 3844 12649 3878
rect 12649 3844 12653 3878
rect 12475 3810 12653 3844
rect 12475 3776 12479 3810
rect 12479 3776 12547 3810
rect 12547 3776 12581 3810
rect 12581 3776 12649 3810
rect 12649 3776 12653 3810
rect 12475 3742 12653 3776
rect 12475 3708 12479 3742
rect 12479 3708 12547 3742
rect 12547 3708 12581 3742
rect 12581 3708 12649 3742
rect 12649 3708 12653 3742
rect 12475 3674 12653 3708
rect 12475 3640 12479 3674
rect 12479 3640 12547 3674
rect 12547 3640 12581 3674
rect 12581 3640 12649 3674
rect 12649 3640 12653 3674
rect 12475 3606 12653 3640
rect 12475 3572 12479 3606
rect 12479 3572 12547 3606
rect 12547 3572 12581 3606
rect 12581 3572 12649 3606
rect 12649 3572 12653 3606
rect 12475 3538 12653 3572
rect 12475 3504 12479 3538
rect 12479 3504 12547 3538
rect 12547 3504 12581 3538
rect 12581 3504 12649 3538
rect 12649 3504 12653 3538
rect 12475 3470 12653 3504
rect 12475 3436 12479 3470
rect 12479 3436 12547 3470
rect 12547 3436 12581 3470
rect 12581 3436 12649 3470
rect 12649 3436 12653 3470
rect 12475 3402 12653 3436
rect 12475 3368 12479 3402
rect 12479 3368 12547 3402
rect 12547 3368 12581 3402
rect 12581 3368 12649 3402
rect 12649 3368 12653 3402
rect 12475 3334 12653 3368
rect 12475 3300 12479 3334
rect 12479 3300 12547 3334
rect 12547 3300 12581 3334
rect 12581 3300 12649 3334
rect 12649 3300 12653 3334
rect 12475 3266 12653 3300
rect 12475 3232 12479 3266
rect 12479 3232 12547 3266
rect 12547 3232 12581 3266
rect 12581 3232 12649 3266
rect 12649 3232 12653 3266
rect 12475 3198 12653 3232
rect 12475 3194 12479 3198
rect 12479 3194 12547 3198
rect 12547 3194 12581 3198
rect 12581 3194 12649 3198
rect 12649 3194 12653 3198
rect 12547 3164 12581 3182
rect 12547 3148 12581 3164
rect 12475 3074 12509 3108
rect 12547 3074 12581 3108
rect 12619 3074 12653 3108
rect 12475 2994 12509 3028
rect 12547 2994 12581 3028
rect 12619 2994 12653 3028
rect 12475 2914 12509 2948
rect 12547 2914 12581 2948
rect 12619 2914 12653 2948
rect 12475 2834 12509 2868
rect 12547 2834 12581 2868
rect 12619 2834 12653 2868
rect 12475 2754 12509 2788
rect 12547 2754 12581 2788
rect 12619 2754 12653 2788
rect 12475 2674 12509 2708
rect 12547 2674 12581 2708
rect 12619 2674 12653 2708
rect 12475 2594 12509 2628
rect 12547 2594 12581 2628
rect 12619 2594 12653 2628
rect 12547 2540 12581 2556
rect 12547 2522 12581 2540
rect 12475 2506 12479 2518
rect 12479 2506 12547 2518
rect 12547 2506 12581 2518
rect 12581 2506 12649 2518
rect 12649 2506 12653 2518
rect 12475 2472 12653 2506
rect 12475 2438 12479 2472
rect 12479 2438 12547 2472
rect 12547 2438 12581 2472
rect 12581 2438 12649 2472
rect 12649 2438 12653 2472
rect 12475 2404 12653 2438
rect 12475 2370 12479 2404
rect 12479 2370 12547 2404
rect 12547 2370 12581 2404
rect 12581 2370 12649 2404
rect 12649 2370 12653 2404
rect 12475 2336 12653 2370
rect 12475 2302 12479 2336
rect 12479 2302 12547 2336
rect 12547 2302 12581 2336
rect 12581 2302 12649 2336
rect 12649 2302 12653 2336
rect 12475 2268 12653 2302
rect 12475 2234 12479 2268
rect 12479 2234 12547 2268
rect 12547 2234 12581 2268
rect 12581 2234 12649 2268
rect 12649 2234 12653 2268
rect 12475 2200 12653 2234
rect 12475 2166 12479 2200
rect 12479 2166 12547 2200
rect 12547 2166 12581 2200
rect 12581 2166 12649 2200
rect 12649 2166 12653 2200
rect 12475 2132 12653 2166
rect 12475 2098 12479 2132
rect 12479 2098 12547 2132
rect 12547 2098 12581 2132
rect 12581 2098 12649 2132
rect 12649 2098 12653 2132
rect 12475 2064 12653 2098
rect 12475 2030 12479 2064
rect 12479 2030 12547 2064
rect 12547 2030 12581 2064
rect 12581 2030 12649 2064
rect 12649 2030 12653 2064
rect 12475 1996 12653 2030
rect 12475 1962 12479 1996
rect 12479 1962 12547 1996
rect 12547 1962 12581 1996
rect 12581 1962 12649 1996
rect 12649 1962 12653 1996
rect 12475 1928 12653 1962
rect 12475 1894 12479 1928
rect 12479 1894 12547 1928
rect 12547 1894 12581 1928
rect 12581 1894 12649 1928
rect 12649 1894 12653 1928
rect 12475 1860 12653 1894
rect 12475 1826 12479 1860
rect 12479 1826 12547 1860
rect 12547 1826 12581 1860
rect 12581 1826 12649 1860
rect 12649 1826 12653 1860
rect 12475 1792 12653 1826
rect 12475 1758 12479 1792
rect 12479 1758 12547 1792
rect 12547 1758 12581 1792
rect 12581 1758 12649 1792
rect 12649 1758 12653 1792
rect 12475 1724 12653 1758
rect 12475 1690 12479 1724
rect 12479 1690 12547 1724
rect 12547 1690 12581 1724
rect 12581 1690 12649 1724
rect 12649 1690 12653 1724
rect 12475 1656 12653 1690
rect 12475 1622 12479 1656
rect 12479 1622 12547 1656
rect 12547 1622 12581 1656
rect 12581 1622 12649 1656
rect 12649 1622 12653 1656
rect 12475 1620 12653 1622
rect 12547 1586 12581 1620
rect 12230 1144 12336 1250
rect 12971 4064 13005 4098
rect 13043 4064 13077 4098
rect 13115 4064 13149 4098
rect 12971 3991 13005 4025
rect 13043 3991 13077 4025
rect 13115 3991 13149 4025
rect 12971 3918 13005 3952
rect 13043 3918 13077 3952
rect 13115 3918 13149 3952
rect 12971 3845 13005 3879
rect 13043 3845 13077 3879
rect 13115 3845 13149 3879
rect 12971 3772 13005 3806
rect 13043 3772 13077 3806
rect 13115 3772 13149 3806
rect 12971 3699 13005 3733
rect 13043 3699 13077 3733
rect 13115 3699 13149 3733
rect 12971 3626 13005 3660
rect 13043 3626 13077 3660
rect 13115 3626 13149 3660
rect 12971 3553 13005 3587
rect 13043 3553 13077 3587
rect 13115 3553 13149 3587
rect 12971 3480 13005 3514
rect 13043 3480 13077 3514
rect 13115 3480 13149 3514
rect 12971 3407 13005 3441
rect 13043 3407 13077 3441
rect 13115 3407 13149 3441
rect 12971 3334 13005 3368
rect 13043 3334 13077 3368
rect 13115 3334 13149 3368
rect 12971 3261 13005 3295
rect 13043 3261 13077 3295
rect 13115 3261 13149 3295
rect 12971 3188 13005 3222
rect 13043 3188 13077 3222
rect 13115 3188 13149 3222
rect 12971 3115 13005 3149
rect 13043 3115 13077 3149
rect 13115 3115 13149 3149
rect 12971 3042 13005 3076
rect 13043 3042 13077 3076
rect 13115 3042 13149 3076
rect 12971 2969 13005 3003
rect 13043 2969 13077 3003
rect 13115 2969 13149 3003
rect 12971 2896 13005 2930
rect 13043 2896 13077 2930
rect 13115 2896 13149 2930
rect 12971 2823 13005 2857
rect 13043 2823 13077 2857
rect 13115 2823 13149 2857
rect 12971 2750 13005 2784
rect 13043 2750 13077 2784
rect 13115 2750 13149 2784
rect 12971 2677 13005 2711
rect 13043 2677 13077 2711
rect 13115 2677 13149 2711
rect 12971 2604 13005 2638
rect 13043 2604 13077 2638
rect 13115 2604 13149 2638
rect 12971 2531 13005 2565
rect 13043 2531 13077 2565
rect 13115 2531 13149 2565
rect 12971 2458 13005 2492
rect 13043 2458 13077 2492
rect 13115 2458 13149 2492
rect 12971 2385 13005 2419
rect 13043 2385 13077 2419
rect 13115 2385 13149 2419
rect 12971 2312 13005 2346
rect 13043 2312 13077 2346
rect 13115 2312 13149 2346
rect 12971 2239 13005 2273
rect 13043 2239 13077 2273
rect 13115 2239 13149 2273
rect 12971 2166 13005 2200
rect 13043 2166 13077 2200
rect 13115 2166 13149 2200
rect 12971 2092 13005 2126
rect 13043 2092 13077 2126
rect 13115 2092 13149 2126
rect 12971 2018 13005 2052
rect 13043 2018 13077 2052
rect 13115 2018 13149 2052
rect 12971 1944 13005 1978
rect 13043 1944 13077 1978
rect 13115 1944 13149 1978
rect 12971 1870 13005 1904
rect 13043 1870 13077 1904
rect 13115 1870 13149 1904
rect 12971 1796 13005 1830
rect 13043 1796 13077 1830
rect 13115 1796 13149 1830
rect 12971 1722 13005 1756
rect 13043 1722 13077 1756
rect 13115 1722 13149 1756
rect 12971 1648 13005 1682
rect 13043 1648 13077 1682
rect 13115 1648 13149 1682
rect 12971 1574 13005 1608
rect 13043 1574 13077 1608
rect 13115 1574 13149 1608
rect 12792 1144 12898 1250
rect 13539 4092 13573 4118
rect 13467 4082 13645 4092
rect 13467 4048 13471 4082
rect 13471 4048 13539 4082
rect 13539 4048 13573 4082
rect 13573 4048 13641 4082
rect 13641 4048 13645 4082
rect 13467 4014 13645 4048
rect 13467 3980 13471 4014
rect 13471 3980 13539 4014
rect 13539 3980 13573 4014
rect 13573 3980 13641 4014
rect 13641 3980 13645 4014
rect 13467 3946 13645 3980
rect 13467 3912 13471 3946
rect 13471 3912 13539 3946
rect 13539 3912 13573 3946
rect 13573 3912 13641 3946
rect 13641 3912 13645 3946
rect 13467 3878 13645 3912
rect 13467 3844 13471 3878
rect 13471 3844 13539 3878
rect 13539 3844 13573 3878
rect 13573 3844 13641 3878
rect 13641 3844 13645 3878
rect 13467 3810 13645 3844
rect 13467 3776 13471 3810
rect 13471 3776 13539 3810
rect 13539 3776 13573 3810
rect 13573 3776 13641 3810
rect 13641 3776 13645 3810
rect 13467 3742 13645 3776
rect 13467 3708 13471 3742
rect 13471 3708 13539 3742
rect 13539 3708 13573 3742
rect 13573 3708 13641 3742
rect 13641 3708 13645 3742
rect 13467 3674 13645 3708
rect 13467 3640 13471 3674
rect 13471 3640 13539 3674
rect 13539 3640 13573 3674
rect 13573 3640 13641 3674
rect 13641 3640 13645 3674
rect 13467 3606 13645 3640
rect 13467 3572 13471 3606
rect 13471 3572 13539 3606
rect 13539 3572 13573 3606
rect 13573 3572 13641 3606
rect 13641 3572 13645 3606
rect 13467 3538 13645 3572
rect 13467 3504 13471 3538
rect 13471 3504 13539 3538
rect 13539 3504 13573 3538
rect 13573 3504 13641 3538
rect 13641 3504 13645 3538
rect 13467 3470 13645 3504
rect 13467 3436 13471 3470
rect 13471 3436 13539 3470
rect 13539 3436 13573 3470
rect 13573 3436 13641 3470
rect 13641 3436 13645 3470
rect 13467 3402 13645 3436
rect 13467 3368 13471 3402
rect 13471 3368 13539 3402
rect 13539 3368 13573 3402
rect 13573 3368 13641 3402
rect 13641 3368 13645 3402
rect 13467 3334 13645 3368
rect 13467 3300 13471 3334
rect 13471 3300 13539 3334
rect 13539 3300 13573 3334
rect 13573 3300 13641 3334
rect 13641 3300 13645 3334
rect 13467 3266 13645 3300
rect 13467 3232 13471 3266
rect 13471 3232 13539 3266
rect 13539 3232 13573 3266
rect 13573 3232 13641 3266
rect 13641 3232 13645 3266
rect 13467 3198 13645 3232
rect 13467 3194 13471 3198
rect 13471 3194 13539 3198
rect 13539 3194 13573 3198
rect 13573 3194 13641 3198
rect 13641 3194 13645 3198
rect 13539 3164 13573 3182
rect 13539 3148 13573 3164
rect 13467 3074 13501 3108
rect 13539 3074 13573 3108
rect 13611 3074 13645 3108
rect 13467 2994 13501 3028
rect 13539 2994 13573 3028
rect 13611 2994 13645 3028
rect 13467 2914 13501 2948
rect 13539 2914 13573 2948
rect 13611 2914 13645 2948
rect 13467 2834 13501 2868
rect 13539 2834 13573 2868
rect 13611 2834 13645 2868
rect 13467 2754 13501 2788
rect 13539 2754 13573 2788
rect 13611 2754 13645 2788
rect 13467 2674 13501 2708
rect 13539 2674 13573 2708
rect 13611 2674 13645 2708
rect 13467 2594 13501 2628
rect 13539 2594 13573 2628
rect 13611 2594 13645 2628
rect 13539 2540 13573 2556
rect 13539 2522 13573 2540
rect 13467 2506 13471 2518
rect 13471 2506 13539 2518
rect 13539 2506 13573 2518
rect 13573 2506 13641 2518
rect 13641 2506 13645 2518
rect 13467 2472 13645 2506
rect 13467 2438 13471 2472
rect 13471 2438 13539 2472
rect 13539 2438 13573 2472
rect 13573 2438 13641 2472
rect 13641 2438 13645 2472
rect 13467 2404 13645 2438
rect 13467 2370 13471 2404
rect 13471 2370 13539 2404
rect 13539 2370 13573 2404
rect 13573 2370 13641 2404
rect 13641 2370 13645 2404
rect 13467 2336 13645 2370
rect 13467 2302 13471 2336
rect 13471 2302 13539 2336
rect 13539 2302 13573 2336
rect 13573 2302 13641 2336
rect 13641 2302 13645 2336
rect 13467 2268 13645 2302
rect 13467 2234 13471 2268
rect 13471 2234 13539 2268
rect 13539 2234 13573 2268
rect 13573 2234 13641 2268
rect 13641 2234 13645 2268
rect 13467 2200 13645 2234
rect 13467 2166 13471 2200
rect 13471 2166 13539 2200
rect 13539 2166 13573 2200
rect 13573 2166 13641 2200
rect 13641 2166 13645 2200
rect 13467 2132 13645 2166
rect 13467 2098 13471 2132
rect 13471 2098 13539 2132
rect 13539 2098 13573 2132
rect 13573 2098 13641 2132
rect 13641 2098 13645 2132
rect 13467 2064 13645 2098
rect 13467 2030 13471 2064
rect 13471 2030 13539 2064
rect 13539 2030 13573 2064
rect 13573 2030 13641 2064
rect 13641 2030 13645 2064
rect 13467 1996 13645 2030
rect 13467 1962 13471 1996
rect 13471 1962 13539 1996
rect 13539 1962 13573 1996
rect 13573 1962 13641 1996
rect 13641 1962 13645 1996
rect 13467 1928 13645 1962
rect 13467 1894 13471 1928
rect 13471 1894 13539 1928
rect 13539 1894 13573 1928
rect 13573 1894 13641 1928
rect 13641 1894 13645 1928
rect 13467 1860 13645 1894
rect 13467 1826 13471 1860
rect 13471 1826 13539 1860
rect 13539 1826 13573 1860
rect 13573 1826 13641 1860
rect 13641 1826 13645 1860
rect 13467 1792 13645 1826
rect 13467 1758 13471 1792
rect 13471 1758 13539 1792
rect 13539 1758 13573 1792
rect 13573 1758 13641 1792
rect 13641 1758 13645 1792
rect 13467 1724 13645 1758
rect 13467 1690 13471 1724
rect 13471 1690 13539 1724
rect 13539 1690 13573 1724
rect 13573 1690 13641 1724
rect 13641 1690 13645 1724
rect 13467 1656 13645 1690
rect 13467 1622 13471 1656
rect 13471 1622 13539 1656
rect 13539 1622 13573 1656
rect 13573 1622 13641 1656
rect 13641 1622 13645 1656
rect 13467 1620 13645 1622
rect 13539 1586 13573 1620
rect 13222 1144 13328 1250
rect 13999 4082 14033 4098
rect 13999 4064 14033 4082
rect 13999 4014 14033 4025
rect 13999 3991 14033 4014
rect 13999 3946 14033 3952
rect 13999 3918 14033 3946
rect 13999 3878 14033 3879
rect 13999 3845 14033 3878
rect 13999 3776 14033 3806
rect 13999 3772 14033 3776
rect 13999 3708 14033 3733
rect 13999 3699 14033 3708
rect 13999 3640 14033 3660
rect 13999 3626 14033 3640
rect 13999 3572 14033 3587
rect 13999 3553 14033 3572
rect 13999 3504 14033 3514
rect 13999 3480 14033 3504
rect 13999 3436 14033 3441
rect 13999 3407 14033 3436
rect 13999 3334 14033 3368
rect 13999 3266 14033 3295
rect 13999 3261 14033 3266
rect 13999 3198 14033 3222
rect 13999 3188 14033 3198
rect 13999 3115 14033 3149
rect 13999 3042 14033 3076
rect 13999 2969 14033 3003
rect 13999 2896 14033 2930
rect 13999 2823 14033 2857
rect 13999 2750 14033 2784
rect 13999 2677 14033 2711
rect 13999 2604 14033 2638
rect 13999 2531 14033 2565
rect 13999 2482 14033 2492
rect 13999 2458 14033 2482
rect 13999 2414 14033 2419
rect 13999 2385 14033 2414
rect 13999 2312 14033 2346
rect 13999 2244 14033 2273
rect 13999 2239 14033 2244
rect 13999 2176 14033 2200
rect 13999 2166 14033 2176
rect 13999 2108 14033 2126
rect 13999 2092 14033 2108
rect 13999 2040 14033 2052
rect 13999 2018 14033 2040
rect 13999 1972 14033 1978
rect 13999 1944 14033 1972
rect 13999 1870 14033 1904
rect 13999 1802 14033 1830
rect 13999 1796 14033 1802
rect 13999 1734 14033 1756
rect 13999 1722 14033 1734
rect 13999 1666 14033 1682
rect 13999 1648 14033 1666
rect 13999 1598 14033 1608
rect 13999 1574 14033 1598
rect 13784 1144 13890 1250
rect 14142 1144 14248 1250
rect 14356 4252 14390 4286
rect 14356 4179 14390 4213
rect 14356 4106 14390 4140
rect 14356 4048 14390 4067
rect 14356 4033 14390 4048
rect 14356 3980 14390 3994
rect 14356 3960 14390 3980
rect 14428 3992 14468 4426
rect 14468 3992 14606 4426
rect 14428 3960 14536 3992
rect 14536 3960 14606 3992
rect 14356 3912 14390 3921
rect 14428 3918 14462 3952
rect 14356 3887 14390 3912
rect 14500 3888 14534 3921
rect 14572 3905 14604 3921
rect 14604 3905 14606 3921
rect 14500 3887 14502 3888
rect 14502 3887 14534 3888
rect 14356 3844 14390 3848
rect 14428 3846 14462 3880
rect 14572 3887 14606 3905
rect 14356 3814 14390 3844
rect 14500 3819 14534 3848
rect 14572 3837 14604 3848
rect 14604 3837 14606 3848
rect 14500 3814 14502 3819
rect 14502 3814 14534 3819
rect 14356 3742 14390 3775
rect 14428 3774 14462 3808
rect 14572 3814 14606 3837
rect 14500 3750 14534 3775
rect 14572 3769 14604 3775
rect 14604 3769 14606 3775
rect 14356 3741 14390 3742
rect 14500 3741 14502 3750
rect 14502 3741 14534 3750
rect 14428 3702 14462 3736
rect 14572 3741 14606 3769
rect 14356 3674 14390 3702
rect 14500 3681 14534 3702
rect 14572 3701 14604 3702
rect 14604 3701 14606 3702
rect 14356 3668 14390 3674
rect 14500 3668 14502 3681
rect 14502 3668 14534 3681
rect 14428 3630 14462 3664
rect 14572 3668 14606 3701
rect 14356 3606 14390 3629
rect 14500 3612 14534 3629
rect 14356 3595 14390 3606
rect 14500 3595 14502 3612
rect 14502 3595 14534 3612
rect 14428 3558 14462 3592
rect 14572 3599 14606 3629
rect 14572 3595 14604 3599
rect 14604 3595 14606 3599
rect 14356 3538 14390 3556
rect 14500 3543 14534 3556
rect 14356 3522 14390 3538
rect 14500 3522 14502 3543
rect 14502 3522 14534 3543
rect 14428 3486 14462 3520
rect 14572 3531 14606 3556
rect 14572 3522 14604 3531
rect 14604 3522 14606 3531
rect 14356 3470 14390 3483
rect 14500 3474 14534 3483
rect 14356 3449 14390 3470
rect 14500 3449 14502 3474
rect 14502 3449 14534 3474
rect 14428 3414 14462 3448
rect 14572 3463 14606 3483
rect 14572 3449 14604 3463
rect 14604 3449 14606 3463
rect 14356 3402 14390 3410
rect 14500 3405 14534 3410
rect 14356 3376 14390 3402
rect 14500 3376 14502 3405
rect 14502 3376 14534 3405
rect 14428 3342 14462 3376
rect 14572 3395 14606 3410
rect 14572 3376 14604 3395
rect 14604 3376 14606 3395
rect 14356 3334 14390 3337
rect 14500 3336 14534 3337
rect 14356 3303 14390 3334
rect 14428 3270 14462 3304
rect 14500 3303 14502 3336
rect 14502 3303 14534 3336
rect 14572 3327 14606 3337
rect 14572 3303 14604 3327
rect 14604 3303 14606 3327
rect 14356 3232 14390 3264
rect 14500 3233 14502 3264
rect 14502 3233 14534 3264
rect 14572 3259 14606 3264
rect 14356 3230 14390 3232
rect 14428 3198 14462 3232
rect 14500 3230 14534 3233
rect 14572 3230 14604 3259
rect 14604 3230 14606 3259
rect 14356 3164 14390 3191
rect 14500 3164 14502 3191
rect 14502 3164 14534 3191
rect 14356 3157 14390 3164
rect 14428 3126 14462 3160
rect 14500 3157 14534 3164
rect 14572 3157 14604 3191
rect 14604 3157 14606 3191
rect 14356 3084 14390 3118
rect 14500 3095 14502 3118
rect 14502 3095 14534 3118
rect 14428 3054 14462 3088
rect 14500 3084 14534 3095
rect 14572 3089 14604 3118
rect 14604 3089 14606 3118
rect 14572 3084 14606 3089
rect 14356 3011 14390 3045
rect 14500 3026 14502 3045
rect 14502 3026 14534 3045
rect 14428 2982 14462 3016
rect 14500 3011 14534 3026
rect 14572 3021 14604 3045
rect 14604 3021 14606 3045
rect 14572 3011 14606 3021
rect 14356 2938 14390 2972
rect 14500 2957 14502 2972
rect 14502 2957 14534 2972
rect 14428 2910 14462 2944
rect 14500 2938 14534 2957
rect 14572 2953 14604 2972
rect 14604 2953 14606 2972
rect 14572 2938 14606 2953
rect 14356 2865 14390 2899
rect 14500 2888 14502 2899
rect 14502 2888 14534 2899
rect 14428 2838 14462 2872
rect 14500 2865 14534 2888
rect 14572 2885 14604 2899
rect 14604 2885 14606 2899
rect 14572 2865 14606 2885
rect 14356 2792 14390 2826
rect 14500 2819 14502 2826
rect 14502 2819 14534 2826
rect 14428 2766 14462 2800
rect 14500 2792 14534 2819
rect 14572 2817 14604 2826
rect 14604 2817 14606 2826
rect 14572 2792 14606 2817
rect 14356 2719 14390 2753
rect 14500 2750 14502 2753
rect 14502 2750 14534 2753
rect 14428 2694 14462 2728
rect 14500 2719 14534 2750
rect 14572 2749 14604 2753
rect 14604 2749 14606 2753
rect 14572 2719 14606 2749
rect 14356 2646 14390 2680
rect 14428 2622 14462 2656
rect 14500 2646 14534 2680
rect 14572 2647 14606 2680
rect 14572 2646 14604 2647
rect 14604 2646 14606 2647
rect 14356 2573 14390 2607
rect 14428 2550 14462 2584
rect 14500 2577 14534 2607
rect 14572 2579 14606 2607
rect 14500 2573 14502 2577
rect 14502 2573 14534 2577
rect 14572 2573 14604 2579
rect 14604 2573 14606 2579
rect 14356 2500 14390 2534
rect 14428 2478 14462 2512
rect 14500 2508 14534 2534
rect 14572 2511 14606 2534
rect 14500 2500 14502 2508
rect 14502 2500 14534 2508
rect 14572 2500 14604 2511
rect 14604 2500 14606 2511
rect 14356 2448 14390 2461
rect 14356 2427 14390 2448
rect 14428 2406 14462 2440
rect 14500 2439 14534 2461
rect 14572 2443 14606 2461
rect 14500 2427 14502 2439
rect 14502 2427 14534 2439
rect 14572 2427 14604 2443
rect 14604 2427 14606 2443
rect 14356 2380 14390 2388
rect 14356 2354 14390 2380
rect 14500 2370 14534 2388
rect 14572 2375 14606 2388
rect 14428 2334 14462 2368
rect 14500 2354 14502 2370
rect 14502 2354 14534 2370
rect 14572 2354 14604 2375
rect 14604 2354 14606 2375
rect 14356 2312 14390 2315
rect 14356 2281 14390 2312
rect 14500 2301 14534 2315
rect 14572 2307 14606 2315
rect 14428 2262 14462 2296
rect 14500 2281 14502 2301
rect 14502 2281 14534 2301
rect 14572 2281 14604 2307
rect 14604 2281 14606 2307
rect 14356 2210 14390 2242
rect 14500 2232 14534 2242
rect 14572 2239 14606 2242
rect 14356 2208 14390 2210
rect 14428 2190 14462 2224
rect 14500 2208 14502 2232
rect 14502 2208 14534 2232
rect 14572 2208 14604 2239
rect 14604 2208 14606 2239
rect 14356 2142 14390 2169
rect 14500 2163 14534 2169
rect 14356 2135 14390 2142
rect 14428 2118 14462 2152
rect 14500 2135 14502 2163
rect 14502 2135 14534 2163
rect 14572 2137 14604 2169
rect 14604 2137 14606 2169
rect 14572 2135 14606 2137
rect 14356 2074 14390 2096
rect 14500 2094 14534 2096
rect 14356 2062 14390 2074
rect 14428 2046 14462 2080
rect 14500 2062 14502 2094
rect 14502 2062 14534 2094
rect 14572 2069 14604 2096
rect 14604 2069 14606 2096
rect 14572 2062 14606 2069
rect 14356 2006 14390 2023
rect 14356 1989 14390 2006
rect 14428 1974 14462 2008
rect 14500 1991 14502 2023
rect 14502 1991 14534 2023
rect 14572 2001 14604 2023
rect 14604 2001 14606 2023
rect 14500 1989 14534 1991
rect 14572 1989 14606 2001
rect 14356 1938 14390 1950
rect 14356 1916 14390 1938
rect 14428 1902 14462 1936
rect 14500 1922 14502 1950
rect 14502 1922 14534 1950
rect 14572 1933 14604 1950
rect 14604 1933 14606 1950
rect 14500 1916 14534 1922
rect 14572 1916 14606 1933
rect 14356 1870 14390 1877
rect 14356 1843 14390 1870
rect 14428 1830 14462 1864
rect 14500 1853 14502 1877
rect 14502 1853 14534 1877
rect 14572 1865 14604 1877
rect 14604 1865 14606 1877
rect 14500 1843 14534 1853
rect 14572 1843 14606 1865
rect 14356 1802 14390 1804
rect 14356 1770 14390 1802
rect 14428 1758 14462 1792
rect 14500 1784 14502 1804
rect 14502 1784 14534 1804
rect 14572 1797 14604 1804
rect 14604 1797 14606 1804
rect 14500 1770 14534 1784
rect 14572 1770 14606 1797
rect 14356 1700 14390 1731
rect 14356 1697 14390 1700
rect 14428 1686 14462 1720
rect 14500 1715 14502 1731
rect 14502 1715 14534 1731
rect 14572 1729 14604 1731
rect 14604 1729 14606 1731
rect 14500 1697 14534 1715
rect 14572 1697 14606 1729
rect 14356 1632 14390 1657
rect 14356 1623 14390 1632
rect 14428 1614 14462 1648
rect 14500 1646 14502 1658
rect 14502 1646 14534 1658
rect 14500 1624 14534 1646
rect 14572 1627 14606 1658
rect 14572 1624 14604 1627
rect 14604 1624 14606 1627
rect 14356 1564 14390 1583
rect 14500 1577 14502 1585
rect 14502 1577 14534 1585
rect 14356 1549 14390 1564
rect 14428 1542 14462 1576
rect 14500 1551 14534 1577
rect 14572 1559 14606 1585
rect 14572 1551 14604 1559
rect 14604 1551 14606 1559
rect 14356 1475 14390 1509
rect 14500 1508 14502 1512
rect 14502 1508 14534 1512
rect 14428 1470 14462 1504
rect 14500 1478 14534 1508
rect 14572 1491 14606 1512
rect 14572 1478 14604 1491
rect 14604 1478 14606 1491
rect 14356 1401 14390 1435
rect 14428 1398 14462 1432
rect 14500 1405 14534 1439
rect 14572 1423 14606 1439
rect 14572 1405 14604 1423
rect 14604 1405 14606 1423
rect 14356 1327 14390 1361
rect 14428 1326 14462 1360
rect 14500 1335 14534 1366
rect 14572 1355 14606 1366
rect 14500 1332 14502 1335
rect 14502 1332 14534 1335
rect 14572 1332 14604 1355
rect 14604 1332 14606 1355
rect 14356 1253 14390 1287
rect 14428 1254 14462 1288
rect 14500 1266 14534 1293
rect 14572 1287 14606 1293
rect 14500 1259 14502 1266
rect 14502 1259 14534 1266
rect 14572 1259 14604 1287
rect 14604 1259 14606 1287
rect 14356 1179 14390 1213
rect 14428 1182 14462 1216
rect 14500 1197 14534 1220
rect 14572 1218 14606 1220
rect 14500 1186 14502 1197
rect 14502 1186 14534 1197
rect 14572 1186 14604 1218
rect 14604 1186 14606 1218
rect 746 883 780 894
rect 14356 1105 14390 1139
rect 14428 1110 14462 1144
rect 14500 1128 14534 1147
rect 14500 1113 14502 1128
rect 14502 1113 14534 1128
rect 14572 1115 14604 1147
rect 14604 1115 14606 1147
rect 14572 1113 14606 1115
rect 14356 1031 14390 1065
rect 14428 1038 14462 1072
rect 14500 1059 14534 1074
rect 14500 1040 14502 1059
rect 14502 1040 14534 1059
rect 14572 1046 14604 1074
rect 14604 1046 14606 1074
rect 14572 1040 14606 1046
rect 14356 957 14390 991
rect 14428 966 14462 1000
rect 14500 990 14534 1001
rect 14500 967 14502 990
rect 14502 967 14534 990
rect 14572 977 14604 1001
rect 14604 977 14606 1001
rect 14572 967 14606 977
rect 14356 883 14390 917
rect 14428 894 14462 928
rect 14500 921 14534 928
rect 14500 894 14502 921
rect 14502 894 14534 921
rect 14572 908 14604 928
rect 14604 908 14606 928
rect 14572 894 14606 908
rect 709 818 736 820
rect 736 818 743 820
rect 782 818 805 820
rect 805 818 816 820
rect 855 818 874 820
rect 874 818 889 820
rect 928 818 943 820
rect 943 818 978 820
rect 978 818 1012 820
rect 1012 818 1047 820
rect 1047 818 1081 820
rect 1081 818 1116 820
rect 1116 818 1150 820
rect 1150 818 1185 820
rect 1185 818 1219 820
rect 1219 818 1254 820
rect 1254 818 1288 820
rect 1288 818 1323 820
rect 1323 818 1357 820
rect 1357 818 1392 820
rect 1392 818 1426 820
rect 1426 818 1461 820
rect 1461 818 1495 820
rect 1495 818 1530 820
rect 1530 818 1564 820
rect 1564 818 1599 820
rect 1599 818 1633 820
rect 1633 818 1668 820
rect 1668 818 1702 820
rect 1702 818 1737 820
rect 1737 818 1771 820
rect 1771 818 1806 820
rect 1806 818 1840 820
rect 1840 818 1875 820
rect 1875 818 1909 820
rect 1909 818 1944 820
rect 1944 818 1978 820
rect 1978 818 2013 820
rect 2013 818 2047 820
rect 2047 818 2082 820
rect 2082 818 2116 820
rect 2116 818 2151 820
rect 2151 818 2185 820
rect 2185 818 2220 820
rect 2220 818 2254 820
rect 2254 818 2289 820
rect 2289 818 2323 820
rect 2323 818 2358 820
rect 2358 818 2392 820
rect 2392 818 2427 820
rect 2427 818 2461 820
rect 2461 818 2496 820
rect 2496 818 2530 820
rect 2530 818 2565 820
rect 2565 818 2599 820
rect 2599 818 2634 820
rect 2634 818 2668 820
rect 2668 818 2703 820
rect 2703 818 2737 820
rect 2737 818 2772 820
rect 709 786 743 818
rect 782 786 816 818
rect 855 786 889 818
rect 928 784 2772 818
rect 928 750 944 784
rect 944 750 979 784
rect 979 750 1013 784
rect 1013 750 1048 784
rect 1048 750 1082 784
rect 1082 750 1117 784
rect 1117 750 1151 784
rect 1151 750 1186 784
rect 1186 750 1220 784
rect 1220 750 1255 784
rect 1255 750 1289 784
rect 1289 750 1324 784
rect 1324 750 1358 784
rect 1358 750 1393 784
rect 1393 750 1427 784
rect 1427 750 1462 784
rect 1462 750 1496 784
rect 1496 750 1531 784
rect 1531 750 1565 784
rect 1565 750 1600 784
rect 1600 750 1634 784
rect 1634 750 1669 784
rect 1669 750 1703 784
rect 1703 750 1738 784
rect 1738 750 1772 784
rect 1772 750 1807 784
rect 1807 750 1841 784
rect 1841 750 1876 784
rect 1876 750 1910 784
rect 1910 750 1945 784
rect 1945 750 1979 784
rect 1979 750 2014 784
rect 2014 750 2048 784
rect 2048 750 2083 784
rect 2083 750 2117 784
rect 2117 750 2152 784
rect 2152 750 2186 784
rect 2186 750 2221 784
rect 2221 750 2255 784
rect 2255 750 2290 784
rect 2290 750 2324 784
rect 2324 750 2359 784
rect 2359 750 2393 784
rect 2393 750 2428 784
rect 2428 750 2462 784
rect 2462 750 2497 784
rect 2497 750 2531 784
rect 2531 750 2566 784
rect 2566 750 2600 784
rect 2600 750 2635 784
rect 2635 750 2669 784
rect 2669 750 2704 784
rect 2704 750 2738 784
rect 2738 750 2772 784
rect 2772 750 14426 820
rect 709 716 743 748
rect 782 716 816 748
rect 855 716 889 748
rect 928 716 4725 750
rect 709 714 723 716
rect 723 714 743 716
rect 782 714 792 716
rect 792 714 816 716
rect 855 714 861 716
rect 861 714 889 716
rect 928 714 930 716
rect 930 714 964 716
rect 964 714 999 716
rect 999 714 1033 716
rect 1033 714 1068 716
rect 1068 714 1102 716
rect 1102 714 1137 716
rect 1137 714 1171 716
rect 1171 714 1206 716
rect 1206 714 1240 716
rect 1240 714 1275 716
rect 1275 714 1309 716
rect 1309 714 1344 716
rect 1344 714 1378 716
rect 1378 714 1413 716
rect 1413 714 1447 716
rect 1447 714 1482 716
rect 1482 714 1516 716
rect 1516 714 1551 716
rect 1551 714 1585 716
rect 1585 714 1620 716
rect 1620 714 1654 716
rect 1654 714 1689 716
rect 1689 714 1723 716
rect 1723 714 1758 716
rect 1758 714 1792 716
rect 1792 714 1827 716
rect 1827 714 1861 716
rect 1861 714 1896 716
rect 1896 714 1930 716
rect 1930 714 1965 716
rect 1965 714 1999 716
rect 1999 714 2034 716
rect 2034 714 2068 716
rect 2068 714 2103 716
rect 2103 714 2137 716
rect 2137 714 2172 716
rect 2172 714 2206 716
rect 2206 714 2241 716
rect 2241 714 2275 716
rect 2275 714 2310 716
rect 2310 714 2344 716
rect 2344 714 2379 716
rect 2379 714 2413 716
rect 2413 714 2448 716
rect 2448 714 2482 716
rect 2482 714 2517 716
rect 2517 714 2551 716
rect 2551 714 2586 716
rect 2586 714 2620 716
rect 2620 714 2655 716
rect 2655 714 2689 716
rect 2689 714 2724 716
rect 2724 714 2758 716
rect 2758 714 2793 716
rect 2793 714 2827 716
rect 2827 714 2862 716
rect 2862 714 2896 716
rect 2896 714 2931 716
rect 2931 714 2965 716
rect 2965 714 3000 716
rect 3000 714 3034 716
rect 3034 714 3069 716
rect 3069 714 3103 716
rect 3103 714 3138 716
rect 3138 714 3172 716
rect 3172 714 3207 716
rect 3207 714 3241 716
rect 3241 714 3276 716
rect 3276 714 3310 716
rect 3310 714 3345 716
rect 3345 714 3379 716
rect 3379 714 3414 716
rect 3414 714 3448 716
rect 3448 714 3483 716
rect 3483 714 3517 716
rect 3517 714 3552 716
rect 3552 714 3586 716
rect 3586 714 3621 716
rect 3621 714 3655 716
rect 3655 714 3690 716
rect 3690 714 3724 716
rect 3724 714 3759 716
rect 3759 714 3793 716
rect 3793 714 3828 716
rect 3828 714 3862 716
rect 3862 714 3897 716
rect 3897 714 3931 716
rect 3931 714 3966 716
rect 3966 714 4000 716
rect 4000 714 4035 716
rect 4035 714 4069 716
rect 4069 714 4104 716
rect 4104 714 4138 716
rect 4138 714 4173 716
rect 4173 714 4207 716
rect 4207 714 4242 716
rect 4242 714 4276 716
rect 4276 714 4311 716
rect 4311 714 4345 716
rect 4345 714 4380 716
rect 4380 714 4414 716
rect 4414 714 4449 716
rect 4449 714 4483 716
rect 4483 714 4518 716
rect 4518 714 4552 716
rect 4552 714 4587 716
rect 4587 714 4621 716
rect 4621 714 4656 716
rect 4656 714 4690 716
rect 4690 714 4725 716
rect 4725 714 14426 750
rect 14832 4655 14866 4670
rect 14907 4657 15085 4695
rect 14832 4636 14840 4655
rect 14840 4636 14866 4655
rect 14907 4623 14915 4657
rect 14915 4623 14949 4657
rect 14949 4623 14983 4657
rect 14983 4623 15017 4657
rect 15017 4623 15051 4657
rect 15051 4623 15085 4657
rect 14832 4587 14866 4598
rect 14832 4564 14840 4587
rect 14840 4564 14866 4587
rect 14907 4585 15085 4623
rect 14907 4551 14915 4585
rect 14915 4551 14949 4585
rect 14949 4551 14983 4585
rect 14983 4551 15017 4585
rect 15017 4551 15051 4585
rect 15051 4551 15085 4585
rect 14832 4519 14866 4526
rect 14832 4492 14840 4519
rect 14840 4492 14866 4519
rect 14907 4513 15085 4551
rect 14907 4479 14915 4513
rect 14915 4479 14949 4513
rect 14949 4479 14983 4513
rect 14983 4479 15017 4513
rect 15017 4479 15051 4513
rect 15051 4479 15085 4513
rect 14832 4451 14866 4454
rect 14832 4420 14840 4451
rect 14840 4420 14866 4451
rect 14907 4441 15085 4479
rect 14907 4407 14915 4441
rect 14915 4407 14949 4441
rect 14949 4407 14983 4441
rect 14983 4407 15017 4441
rect 15017 4407 15051 4441
rect 15051 4407 15085 4441
rect 14832 4349 14840 4382
rect 14840 4349 14866 4382
rect 14907 4369 15085 4407
rect 14907 4368 14983 4369
rect 14832 4348 14866 4349
rect 14907 4334 14915 4368
rect 14915 4334 14949 4368
rect 14949 4335 14983 4368
rect 14983 4335 15017 4369
rect 15017 4335 15051 4369
rect 15051 4335 15085 4369
rect 14949 4334 15085 4335
rect 14832 4281 14840 4310
rect 14840 4281 14866 4310
rect 14907 4297 15085 4334
rect 14907 4295 14983 4297
rect 14832 4276 14866 4281
rect 14907 4261 14915 4295
rect 14915 4261 14949 4295
rect 14949 4263 14983 4295
rect 14983 4263 15017 4297
rect 15017 4263 15051 4297
rect 15051 4263 15085 4297
rect 14949 4261 15085 4263
rect 14832 4213 14840 4238
rect 14840 4213 14866 4238
rect 14907 4225 15085 4261
rect 14907 4222 14983 4225
rect 14832 4204 14866 4213
rect 14907 4188 14915 4222
rect 14915 4188 14949 4222
rect 14949 4191 14983 4222
rect 14983 4191 15017 4225
rect 15017 4191 15051 4225
rect 15051 4191 15085 4225
rect 14949 4188 15085 4191
rect 14832 4145 14840 4166
rect 14840 4145 14866 4166
rect 14907 4153 15085 4188
rect 14907 4149 14983 4153
rect 14832 4132 14866 4145
rect 14907 4115 14915 4149
rect 14915 4115 14949 4149
rect 14949 4119 14983 4149
rect 14983 4119 15017 4153
rect 15017 4119 15051 4153
rect 15051 4119 15085 4153
rect 14949 4115 15085 4119
rect 14832 4077 14840 4094
rect 14840 4077 14866 4094
rect 14907 4081 15085 4115
rect 14832 4060 14866 4077
rect 14907 4076 14983 4081
rect 14832 4009 14840 4022
rect 14840 4009 14866 4022
rect 14907 4042 14915 4076
rect 14915 4042 14949 4076
rect 14949 4047 14983 4076
rect 14983 4047 15017 4081
rect 15017 4047 15051 4081
rect 15051 4047 15085 4081
rect 14949 4042 15085 4047
rect 14907 4009 15085 4042
rect 14832 3988 14866 4009
rect 14907 4008 15051 4009
rect 14907 4003 14983 4008
rect 14832 3941 14840 3950
rect 14840 3941 14866 3950
rect 14907 3969 14915 4003
rect 14915 3969 14949 4003
rect 14949 3974 14983 4003
rect 14983 3974 15017 4008
rect 15017 3975 15051 4008
rect 15051 3975 15085 4009
rect 15017 3974 15085 3975
rect 14949 3969 15085 3974
rect 14832 3916 14866 3941
rect 14907 3937 15085 3969
rect 14907 3935 15051 3937
rect 14907 3930 14983 3935
rect 14832 3873 14840 3878
rect 14840 3873 14866 3878
rect 14907 3896 14915 3930
rect 14915 3896 14949 3930
rect 14949 3901 14983 3930
rect 14983 3901 15017 3935
rect 15017 3903 15051 3935
rect 15051 3903 15085 3937
rect 15017 3901 15085 3903
rect 14949 3896 15085 3901
rect 14832 3844 14866 3873
rect 14907 3865 15085 3896
rect 14907 3862 15051 3865
rect 14907 3857 14983 3862
rect 14832 3805 14840 3806
rect 14840 3805 14866 3806
rect 14907 3823 14915 3857
rect 14915 3823 14949 3857
rect 14949 3828 14983 3857
rect 14983 3828 15017 3862
rect 15017 3831 15051 3862
rect 15051 3831 15085 3865
rect 15017 3828 15085 3831
rect 14949 3823 15085 3828
rect 14832 3772 14866 3805
rect 14907 3793 15085 3823
rect 14907 3789 15051 3793
rect 14907 3784 14983 3789
rect 14907 3750 14915 3784
rect 14915 3750 14949 3784
rect 14949 3755 14983 3784
rect 14983 3755 15017 3789
rect 15017 3759 15051 3789
rect 15051 3759 15085 3793
rect 15017 3755 15085 3759
rect 14949 3750 15085 3755
rect 14832 3703 14866 3734
rect 14907 3721 15085 3750
rect 14907 3716 15051 3721
rect 14907 3711 14983 3716
rect 14832 3700 14840 3703
rect 14840 3700 14866 3703
rect 14907 3677 14915 3711
rect 14915 3677 14949 3711
rect 14949 3682 14983 3711
rect 14983 3682 15017 3716
rect 15017 3687 15051 3716
rect 15051 3687 15085 3721
rect 15017 3682 15085 3687
rect 14949 3677 15085 3682
rect 14832 3635 14866 3662
rect 14907 3649 15085 3677
rect 14907 3643 15051 3649
rect 14907 3638 14983 3643
rect 14832 3628 14840 3635
rect 14840 3628 14866 3635
rect 14907 3604 14915 3638
rect 14915 3604 14949 3638
rect 14949 3609 14983 3638
rect 14983 3609 15017 3643
rect 15017 3615 15051 3643
rect 15051 3615 15085 3649
rect 15017 3609 15085 3615
rect 14949 3604 15085 3609
rect 14832 3567 14866 3590
rect 14907 3577 15085 3604
rect 14907 3570 15051 3577
rect 14832 3556 14840 3567
rect 14840 3556 14866 3567
rect 14907 3565 14983 3570
rect 14907 3531 14915 3565
rect 14915 3531 14949 3565
rect 14949 3536 14983 3565
rect 14983 3536 15017 3570
rect 15017 3543 15051 3570
rect 15051 3543 15085 3577
rect 15017 3536 15085 3543
rect 14949 3531 15085 3536
rect 14832 3499 14866 3518
rect 14907 3505 15085 3531
rect 14832 3484 14840 3499
rect 14840 3484 14866 3499
rect 14907 3497 15051 3505
rect 14907 3492 14983 3497
rect 14907 3458 14915 3492
rect 14915 3458 14949 3492
rect 14949 3463 14983 3492
rect 14983 3463 15017 3497
rect 15017 3471 15051 3497
rect 15051 3471 15085 3505
rect 15017 3463 15085 3471
rect 14949 3458 15085 3463
rect 14832 3431 14866 3446
rect 14907 3433 15085 3458
rect 14832 3412 14840 3431
rect 14840 3412 14866 3431
rect 14907 3424 15051 3433
rect 14907 3419 14983 3424
rect 14907 3385 14915 3419
rect 14915 3385 14949 3419
rect 14949 3390 14983 3419
rect 14983 3390 15017 3424
rect 15017 3399 15051 3424
rect 15051 3399 15085 3433
rect 15017 3390 15085 3399
rect 14949 3385 15085 3390
rect 14832 3363 14866 3374
rect 14832 3340 14840 3363
rect 14840 3340 14866 3363
rect 14907 3361 15085 3385
rect 14907 3351 15051 3361
rect 14907 3346 14983 3351
rect 14907 3312 14915 3346
rect 14915 3312 14949 3346
rect 14949 3317 14983 3346
rect 14983 3317 15017 3351
rect 15017 3327 15051 3351
rect 15051 3327 15085 3361
rect 15017 3317 15085 3327
rect 14949 3312 15085 3317
rect 14832 3295 14866 3302
rect 14832 3268 14840 3295
rect 14840 3268 14866 3295
rect 14907 3289 15085 3312
rect 14907 3278 15051 3289
rect 14907 3273 14983 3278
rect 14907 3239 14915 3273
rect 14915 3239 14949 3273
rect 14949 3244 14983 3273
rect 14983 3244 15017 3278
rect 15017 3255 15051 3278
rect 15051 3255 15085 3289
rect 15017 3244 15085 3255
rect 14949 3239 15085 3244
rect 14832 3227 14866 3230
rect 14832 3196 14840 3227
rect 14840 3196 14866 3227
rect 14907 3217 15085 3239
rect 14907 3205 15051 3217
rect 14907 3200 14983 3205
rect 14907 3166 14915 3200
rect 14915 3166 14949 3200
rect 14949 3171 14983 3200
rect 14983 3171 15017 3205
rect 15017 3183 15051 3205
rect 15051 3183 15085 3217
rect 15017 3171 15085 3183
rect 14949 3166 15085 3171
rect 14832 3125 14840 3158
rect 14840 3125 14866 3158
rect 14907 3145 15085 3166
rect 14907 3132 15051 3145
rect 14907 3127 14983 3132
rect 14832 3124 14866 3125
rect 14907 3093 14915 3127
rect 14915 3093 14949 3127
rect 14949 3098 14983 3127
rect 14983 3098 15017 3132
rect 15017 3111 15051 3132
rect 15051 3111 15085 3145
rect 15017 3098 15085 3111
rect 14949 3093 15085 3098
rect 14832 3057 14840 3086
rect 14840 3057 14866 3086
rect 14907 3073 15085 3093
rect 14907 3059 15051 3073
rect 14832 3052 14866 3057
rect 14907 3054 14983 3059
rect 14832 2989 14840 3014
rect 14840 2989 14866 3014
rect 14907 3020 14915 3054
rect 14915 3020 14949 3054
rect 14949 3025 14983 3054
rect 14983 3025 15017 3059
rect 15017 3039 15051 3059
rect 15051 3039 15085 3073
rect 15017 3025 15085 3039
rect 14949 3020 15085 3025
rect 14907 3001 15085 3020
rect 14832 2980 14866 2989
rect 14907 2986 15051 3001
rect 14907 2981 14983 2986
rect 14832 2921 14840 2942
rect 14840 2921 14866 2942
rect 14907 2947 14915 2981
rect 14915 2947 14949 2981
rect 14949 2952 14983 2981
rect 14983 2952 15017 2986
rect 15017 2967 15051 2986
rect 15051 2967 15085 3001
rect 15017 2952 15085 2967
rect 14949 2947 15085 2952
rect 14907 2929 15085 2947
rect 14832 2908 14866 2921
rect 14907 2913 15051 2929
rect 14907 2908 14983 2913
rect 14832 2853 14840 2870
rect 14840 2853 14866 2870
rect 14907 2874 14915 2908
rect 14915 2874 14949 2908
rect 14949 2879 14983 2908
rect 14983 2879 15017 2913
rect 15017 2895 15051 2913
rect 15051 2895 15085 2929
rect 15017 2879 15085 2895
rect 14949 2874 15085 2879
rect 14907 2857 15085 2874
rect 14832 2836 14866 2853
rect 14907 2840 15051 2857
rect 14907 2835 14983 2840
rect 14832 2785 14840 2798
rect 14840 2785 14866 2798
rect 14907 2801 14915 2835
rect 14915 2801 14949 2835
rect 14949 2806 14983 2835
rect 14983 2806 15017 2840
rect 15017 2823 15051 2840
rect 15051 2823 15085 2857
rect 15017 2806 15085 2823
rect 14949 2801 15085 2806
rect 14907 2785 15085 2801
rect 14832 2764 14866 2785
rect 14907 2767 15051 2785
rect 14907 2762 14983 2767
rect 14832 2717 14840 2726
rect 14840 2717 14866 2726
rect 14907 2728 14915 2762
rect 14915 2728 14949 2762
rect 14949 2733 14983 2762
rect 14983 2733 15017 2767
rect 15017 2751 15051 2767
rect 15051 2751 15085 2785
rect 15017 2733 15085 2751
rect 14949 2728 15085 2733
rect 14832 2692 14866 2717
rect 14907 2713 15085 2728
rect 14907 2694 15051 2713
rect 14907 2689 14983 2694
rect 14832 2649 14840 2654
rect 14840 2649 14866 2654
rect 14907 2655 14915 2689
rect 14915 2655 14949 2689
rect 14949 2660 14983 2689
rect 14983 2660 15017 2694
rect 15017 2679 15051 2694
rect 15051 2679 15085 2713
rect 15017 2660 15085 2679
rect 14949 2655 15085 2660
rect 14832 2620 14866 2649
rect 14907 2641 15085 2655
rect 14907 2621 15051 2641
rect 14907 2616 14983 2621
rect 14832 2581 14840 2582
rect 14840 2581 14866 2582
rect 14907 2582 14915 2616
rect 14915 2582 14949 2616
rect 14949 2587 14983 2616
rect 14983 2587 15017 2621
rect 15017 2607 15051 2621
rect 15051 2607 15085 2641
rect 15017 2587 15085 2607
rect 14949 2582 15085 2587
rect 14832 2548 14866 2581
rect 14907 2569 15085 2582
rect 14907 2548 15051 2569
rect 14907 2543 14983 2548
rect 14832 2479 14866 2510
rect 14907 2509 14915 2543
rect 14915 2509 14949 2543
rect 14949 2514 14983 2543
rect 14983 2514 15017 2548
rect 15017 2535 15051 2548
rect 15051 2535 15085 2569
rect 15017 2514 15085 2535
rect 14949 2509 15085 2514
rect 14907 2497 15085 2509
rect 14832 2476 14840 2479
rect 14840 2476 14866 2479
rect 14907 2475 15051 2497
rect 14907 2470 14983 2475
rect 14832 2411 14866 2438
rect 14907 2436 14915 2470
rect 14915 2436 14949 2470
rect 14949 2441 14983 2470
rect 14983 2441 15017 2475
rect 15017 2463 15051 2475
rect 15051 2463 15085 2497
rect 15017 2441 15085 2463
rect 14949 2436 15085 2441
rect 14907 2425 15085 2436
rect 14832 2404 14840 2411
rect 14840 2404 14866 2411
rect 14907 2402 15051 2425
rect 14907 2397 14983 2402
rect 14832 2343 14866 2366
rect 14907 2363 14915 2397
rect 14915 2363 14949 2397
rect 14949 2368 14983 2397
rect 14983 2368 15017 2402
rect 15017 2391 15051 2402
rect 15051 2391 15085 2425
rect 15017 2368 15085 2391
rect 14949 2363 15085 2368
rect 14907 2353 15085 2363
rect 14832 2332 14840 2343
rect 14840 2332 14866 2343
rect 14907 2329 15051 2353
rect 14907 2324 14983 2329
rect 14832 2275 14866 2294
rect 14907 2290 14915 2324
rect 14915 2290 14949 2324
rect 14949 2295 14983 2324
rect 14983 2295 15017 2329
rect 15017 2319 15051 2329
rect 15051 2319 15085 2353
rect 15017 2295 15085 2319
rect 14949 2290 15085 2295
rect 14907 2280 15085 2290
rect 14832 2260 14840 2275
rect 14840 2260 14866 2275
rect 14907 2256 15051 2280
rect 14907 2251 14983 2256
rect 14832 2207 14866 2222
rect 14907 2217 14915 2251
rect 14915 2217 14949 2251
rect 14949 2222 14983 2251
rect 14983 2222 15017 2256
rect 15017 2246 15051 2256
rect 15051 2246 15085 2280
rect 15017 2222 15085 2246
rect 14949 2217 15085 2222
rect 14907 2207 15085 2217
rect 14832 2188 14840 2207
rect 14840 2188 14866 2207
rect 14907 2183 15051 2207
rect 14907 2178 14983 2183
rect 14832 2139 14866 2150
rect 14907 2144 14915 2178
rect 14915 2144 14949 2178
rect 14949 2149 14983 2178
rect 14983 2149 15017 2183
rect 15017 2173 15051 2183
rect 15051 2173 15085 2207
rect 15017 2149 15085 2173
rect 14949 2144 15085 2149
rect 14832 2116 14840 2139
rect 14840 2116 14866 2139
rect 14907 2134 15085 2144
rect 14907 2110 15051 2134
rect 14907 2105 14983 2110
rect 14832 2071 14866 2078
rect 14907 2071 14915 2105
rect 14915 2071 14949 2105
rect 14949 2076 14983 2105
rect 14983 2076 15017 2110
rect 15017 2100 15051 2110
rect 15051 2100 15085 2134
rect 15017 2076 15085 2100
rect 14949 2071 15085 2076
rect 14832 2044 14840 2071
rect 14840 2044 14866 2071
rect 14907 2061 15085 2071
rect 14907 2037 15051 2061
rect 14907 2032 14983 2037
rect 14832 2003 14866 2006
rect 14832 1972 14840 2003
rect 14840 1972 14866 2003
rect 14907 1998 14915 2032
rect 14915 1998 14949 2032
rect 14949 2003 14983 2032
rect 14983 2003 15017 2037
rect 15017 2027 15051 2037
rect 15051 2027 15085 2061
rect 15017 2003 15085 2027
rect 14949 1998 15085 2003
rect 14907 1988 15085 1998
rect 14907 1964 15051 1988
rect 14907 1959 14983 1964
rect 14832 1901 14840 1934
rect 14840 1901 14866 1934
rect 14907 1925 14915 1959
rect 14915 1925 14949 1959
rect 14949 1930 14983 1959
rect 14983 1930 15017 1964
rect 15017 1954 15051 1964
rect 15051 1954 15085 1988
rect 15017 1930 15085 1954
rect 14949 1925 15085 1930
rect 14907 1915 15085 1925
rect 14832 1900 14866 1901
rect 14907 1891 15051 1915
rect 14907 1886 14983 1891
rect 14832 1833 14840 1862
rect 14840 1833 14866 1862
rect 14907 1852 14915 1886
rect 14915 1852 14949 1886
rect 14949 1857 14983 1886
rect 14983 1857 15017 1891
rect 15017 1881 15051 1891
rect 15051 1881 15085 1915
rect 15017 1857 15085 1881
rect 14949 1852 15085 1857
rect 14907 1842 15085 1852
rect 14832 1828 14866 1833
rect 14907 1818 15051 1842
rect 14907 1813 14983 1818
rect 14832 1765 14840 1790
rect 14840 1765 14866 1790
rect 14907 1779 14915 1813
rect 14915 1779 14949 1813
rect 14949 1784 14983 1813
rect 14983 1784 15017 1818
rect 15017 1808 15051 1818
rect 15051 1808 15085 1842
rect 15017 1784 15085 1808
rect 14949 1779 15085 1784
rect 14907 1769 15085 1779
rect 14832 1756 14866 1765
rect 14907 1745 15051 1769
rect 14907 1740 14983 1745
rect 14832 1697 14840 1718
rect 14840 1697 14866 1718
rect 14907 1706 14915 1740
rect 14915 1706 14949 1740
rect 14949 1711 14983 1740
rect 14983 1711 15017 1745
rect 15017 1735 15051 1745
rect 15051 1735 15085 1769
rect 15017 1711 15085 1735
rect 14949 1706 15085 1711
rect 14832 1684 14866 1697
rect 14907 1696 15085 1706
rect 14907 1672 15051 1696
rect 14907 1667 14983 1672
rect 14832 1629 14840 1646
rect 14840 1629 14866 1646
rect 14907 1633 14915 1667
rect 14915 1633 14949 1667
rect 14949 1638 14983 1667
rect 14983 1638 15017 1672
rect 15017 1662 15051 1672
rect 15051 1662 15085 1696
rect 15017 1638 15085 1662
rect 14949 1633 15085 1638
rect 14832 1612 14866 1629
rect 14907 1623 15085 1633
rect 14907 1599 15051 1623
rect 14832 1561 14840 1574
rect 14840 1561 14866 1574
rect 14907 1594 14983 1599
rect 14832 1540 14866 1561
rect 14907 1560 14915 1594
rect 14915 1560 14949 1594
rect 14949 1565 14983 1594
rect 14983 1565 15017 1599
rect 15017 1589 15051 1599
rect 15051 1589 15085 1623
rect 15017 1565 15085 1589
rect 14949 1560 15085 1565
rect 14907 1550 15085 1560
rect 14832 1493 14840 1502
rect 14840 1493 14866 1502
rect 14907 1526 15051 1550
rect 14907 1521 14983 1526
rect 14832 1468 14866 1493
rect 14907 1487 14915 1521
rect 14915 1487 14949 1521
rect 14949 1492 14983 1521
rect 14983 1492 15017 1526
rect 15017 1516 15051 1526
rect 15051 1516 15085 1550
rect 15017 1492 15085 1516
rect 14949 1487 15085 1492
rect 14907 1477 15085 1487
rect 14832 1425 14840 1429
rect 14840 1425 14866 1429
rect 14907 1453 15051 1477
rect 14907 1448 14983 1453
rect 14832 1395 14866 1425
rect 14907 1414 14915 1448
rect 14915 1414 14949 1448
rect 14949 1419 14983 1448
rect 14983 1419 15017 1453
rect 15017 1443 15051 1453
rect 15051 1443 15085 1477
rect 15017 1419 15085 1443
rect 14949 1414 15085 1419
rect 14907 1404 15085 1414
rect 14907 1380 15051 1404
rect 14907 1375 14983 1380
rect 14832 1323 14866 1356
rect 14907 1341 14915 1375
rect 14915 1341 14949 1375
rect 14949 1346 14983 1375
rect 14983 1346 15017 1380
rect 15017 1370 15051 1380
rect 15051 1370 15085 1404
rect 15017 1346 15085 1370
rect 14949 1341 15085 1346
rect 14907 1331 15085 1341
rect 14832 1322 14840 1323
rect 14840 1322 14866 1323
rect 14907 1307 15051 1331
rect 14907 1302 14983 1307
rect 14832 1255 14866 1283
rect 14907 1268 14915 1302
rect 14915 1268 14949 1302
rect 14949 1273 14983 1302
rect 14983 1273 15017 1307
rect 15017 1297 15051 1307
rect 15051 1297 15085 1331
rect 15017 1273 15085 1297
rect 14949 1268 15085 1273
rect 14907 1258 15085 1268
rect 14832 1249 14840 1255
rect 14840 1249 14866 1255
rect 14907 1234 15051 1258
rect 14907 1229 14983 1234
rect 14832 1187 14866 1210
rect 14907 1195 14915 1229
rect 14915 1195 14949 1229
rect 14949 1200 14983 1229
rect 14983 1200 15017 1234
rect 15017 1224 15051 1234
rect 15051 1224 15085 1258
rect 15017 1200 15085 1224
rect 14949 1195 15085 1200
rect 14832 1176 14840 1187
rect 14840 1176 14866 1187
rect 14907 1185 15085 1195
rect 14907 1161 15051 1185
rect 14907 1156 14983 1161
rect 14832 1119 14866 1137
rect 14907 1122 14915 1156
rect 14915 1122 14949 1156
rect 14949 1127 14983 1156
rect 14983 1127 15017 1161
rect 15017 1151 15051 1161
rect 15051 1151 15085 1185
rect 15017 1127 15085 1151
rect 14949 1122 15085 1127
rect 14832 1103 14840 1119
rect 14840 1103 14866 1119
rect 14907 1112 15085 1122
rect 14907 1088 15051 1112
rect 14907 1083 14983 1088
rect 14832 1051 14866 1064
rect 14832 1030 14840 1051
rect 14840 1030 14866 1051
rect 14907 1049 14915 1083
rect 14915 1049 14949 1083
rect 14949 1054 14983 1083
rect 14983 1054 15017 1088
rect 15017 1078 15051 1088
rect 15051 1078 15085 1112
rect 15017 1054 15085 1078
rect 14949 1049 15085 1054
rect 14907 1039 15085 1049
rect 14907 1015 15051 1039
rect 14907 1010 14983 1015
rect 14832 983 14866 991
rect 14832 957 14840 983
rect 14840 957 14866 983
rect 14907 976 14915 1010
rect 14915 976 14949 1010
rect 14949 981 14983 1010
rect 14983 981 15017 1015
rect 15017 1005 15051 1015
rect 15051 1005 15085 1039
rect 15017 981 15085 1005
rect 14949 976 15085 981
rect 14907 966 15085 976
rect 14907 942 15051 966
rect 14907 937 14983 942
rect 14832 915 14866 918
rect 14832 884 14840 915
rect 14840 884 14866 915
rect 14907 903 14915 937
rect 14915 903 14949 937
rect 14949 908 14983 937
rect 14983 908 15017 942
rect 15017 932 15051 942
rect 15051 932 15085 966
rect 15017 908 15085 932
rect 14949 903 15085 908
rect 14907 893 15085 903
rect 14907 869 15051 893
rect 14907 864 14983 869
rect 14832 813 14840 845
rect 14840 813 14866 845
rect 14907 830 14915 864
rect 14915 830 14949 864
rect 14949 835 14983 864
rect 14983 835 15017 869
rect 15017 859 15051 869
rect 15051 859 15085 893
rect 15017 835 15085 859
rect 14949 830 15085 835
rect 14907 820 15085 830
rect 14832 811 14866 813
rect 14907 796 15051 820
rect 14907 791 14983 796
rect 14832 745 14840 772
rect 14840 745 14866 772
rect 14907 757 14915 791
rect 14915 757 14949 791
rect 14949 762 14983 791
rect 14983 762 15017 796
rect 15017 786 15051 796
rect 15051 786 15085 820
rect 15017 762 15085 786
rect 14949 757 15085 762
rect 14907 747 15085 757
rect 14832 738 14866 745
rect 14907 723 15051 747
rect 14907 718 14983 723
rect 51 576 85 610
rect 85 576 119 610
rect 119 576 153 610
rect 153 576 187 610
rect 187 576 221 610
rect 221 576 229 610
rect 269 609 296 641
rect 296 609 303 641
rect 269 607 303 609
rect 51 538 229 576
rect 269 541 296 567
rect 296 541 303 567
rect 51 504 85 538
rect 85 504 119 538
rect 119 504 153 538
rect 153 504 187 538
rect 187 504 221 538
rect 221 504 229 538
rect 269 533 303 541
rect 14832 677 14840 699
rect 14840 677 14866 699
rect 14907 684 14915 718
rect 14915 684 14949 718
rect 14949 689 14983 718
rect 14983 689 15017 723
rect 15017 713 15051 723
rect 15051 713 15085 747
rect 15017 689 15085 713
rect 14949 684 15085 689
rect 14832 665 14866 677
rect 14907 674 15085 684
rect 14907 650 15051 674
rect 14907 645 14983 650
rect 14832 609 14840 626
rect 14840 609 14866 626
rect 14907 611 14915 645
rect 14915 611 14949 645
rect 14949 616 14983 645
rect 14983 616 15017 650
rect 15017 640 15051 650
rect 15051 640 15085 674
rect 15017 616 15085 640
rect 14949 611 15085 616
rect 14832 592 14866 609
rect 14907 601 15085 611
rect 14907 577 15051 601
rect 14832 541 14840 553
rect 14840 541 14866 553
rect 14907 572 14983 577
rect 14832 519 14866 541
rect 14907 538 14915 572
rect 14915 538 14949 572
rect 14949 543 14983 572
rect 14983 543 15017 577
rect 15017 567 15051 577
rect 15051 567 15085 601
rect 15017 543 15085 567
rect 14949 538 15085 543
rect 14907 528 15085 538
rect 51 466 229 504
rect 14907 504 15051 528
rect 14907 499 14983 504
rect 51 432 85 466
rect 85 432 119 466
rect 119 432 153 466
rect 153 432 187 466
rect 187 432 221 466
rect 221 432 229 466
rect 343 465 375 497
rect 375 465 377 497
rect 419 465 448 497
rect 448 465 453 497
rect 495 465 521 497
rect 521 465 529 497
rect 571 465 594 497
rect 594 465 605 497
rect 648 465 667 497
rect 667 465 682 497
rect 14465 465 14483 481
rect 14483 465 14499 481
rect 14539 465 14555 481
rect 14555 465 14573 481
rect 14613 465 14627 481
rect 14627 465 14647 481
rect 14686 465 14699 481
rect 14699 465 14720 481
rect 14759 465 14771 481
rect 14771 465 14793 481
rect 14907 465 14915 499
rect 14915 465 14949 499
rect 14949 470 14983 499
rect 14983 470 15017 504
rect 15017 494 15051 504
rect 15051 494 15085 528
rect 15017 470 15085 494
rect 14949 465 15085 470
rect 343 463 377 465
rect 419 463 453 465
rect 495 463 529 465
rect 571 463 605 465
rect 648 463 682 465
rect 14465 447 14499 465
rect 14539 447 14573 465
rect 14613 447 14647 465
rect 14686 447 14720 465
rect 14759 447 14793 465
rect 14907 455 15085 465
rect 51 394 229 432
rect 14907 431 15051 455
rect 14907 397 14911 431
rect 14911 397 14945 431
rect 14945 397 14983 431
rect 14983 397 15017 431
rect 15017 421 15051 431
rect 15051 421 15085 455
rect 15017 397 15085 421
rect 51 360 85 394
rect 85 360 119 394
rect 119 360 153 394
rect 153 360 187 394
rect 187 360 221 394
rect 221 360 229 394
rect 14907 382 15085 397
rect 361 363 395 375
rect 434 363 468 375
rect 507 363 541 375
rect 580 363 614 375
rect 653 363 687 375
rect 726 363 760 375
rect 799 363 833 375
rect 872 363 906 375
rect 945 363 979 375
rect 1018 363 1052 375
rect 1091 363 1125 375
rect 1164 363 1198 375
rect 1237 363 1271 375
rect 1310 363 1344 375
rect 1383 363 1417 375
rect 1456 363 1490 375
rect 1529 363 1563 375
rect 1602 363 1636 375
rect 1675 363 1709 375
rect 1748 363 1782 375
rect 1821 363 1855 375
rect 1894 363 1928 375
rect 1967 363 2001 375
rect 2040 363 2074 375
rect 2113 363 2147 375
rect 2186 363 2220 375
rect 2259 363 2293 375
rect 2332 363 2366 375
rect 2405 363 2439 375
rect 2478 363 2512 375
rect 2551 363 2585 375
rect 2624 363 2658 375
rect 2697 363 2731 375
rect 2770 363 2804 375
rect 2843 363 2877 375
rect 2916 363 2950 375
rect 2989 363 3023 375
rect 3062 363 3096 375
rect 3135 363 3169 375
rect 3208 363 3242 375
rect 3281 363 3315 375
rect 3354 363 3388 375
rect 3427 363 3461 375
rect 3500 363 3534 375
rect 3573 363 3607 375
rect 3646 363 3680 375
rect 3719 363 3753 375
rect 3792 363 3826 375
rect 3865 363 3899 375
rect 3938 363 3972 375
rect 4011 363 4045 375
rect 4084 363 4118 375
rect 4157 363 4191 375
rect 4229 363 4263 375
rect 4301 363 4335 375
rect 4373 363 4407 375
rect 4445 363 4479 375
rect 4517 363 4551 375
rect 4589 363 4623 375
rect 4661 363 4695 375
rect 4733 363 4767 375
rect 4805 363 4839 375
rect 4877 363 4911 375
rect 4949 363 4983 375
rect 5021 363 5055 375
rect 5093 363 5127 375
rect 5165 363 5199 375
rect 5237 363 5271 375
rect 5309 363 5343 375
rect 5381 363 5415 375
rect 5453 363 5487 375
rect 5525 363 5559 375
rect 5597 363 5631 375
rect 5669 363 5703 375
rect 5741 363 5775 375
rect 5813 363 5847 375
rect 5885 363 5919 375
rect 5957 363 5991 375
rect 6029 363 6063 375
rect 6101 363 6135 375
rect 6173 363 6207 375
rect 6245 363 6279 375
rect 6317 363 6351 375
rect 6389 363 6423 375
rect 6461 363 6495 375
rect 6533 363 6567 375
rect 6605 363 6639 375
rect 6677 363 6711 375
rect 6749 363 6783 375
rect 6821 363 6855 375
rect 6893 363 6927 375
rect 6965 363 6999 375
rect 7037 363 7071 375
rect 7109 363 7143 375
rect 7181 363 7215 375
rect 7253 363 7287 375
rect 7325 363 7359 375
rect 7397 363 7431 375
rect 7469 363 7503 375
rect 7541 363 7575 375
rect 7613 363 7647 375
rect 7685 363 7719 375
rect 7757 363 7791 375
rect 7829 363 7863 375
rect 7901 363 7935 375
rect 7973 363 8007 375
rect 8045 363 8079 375
rect 8117 363 8151 375
rect 8189 363 8223 375
rect 8261 363 8295 375
rect 8333 363 8367 375
rect 8405 363 8439 375
rect 8477 363 8511 375
rect 8549 363 8583 375
rect 8621 363 8655 375
rect 8693 363 8727 375
rect 8765 363 8799 375
rect 8837 363 8871 375
rect 8909 363 8943 375
rect 8981 363 9015 375
rect 9053 363 9087 375
rect 9125 363 9159 375
rect 9197 363 9231 375
rect 9269 363 9303 375
rect 9341 363 9375 375
rect 9413 363 9447 375
rect 9485 363 9519 375
rect 9557 363 9591 375
rect 9629 363 9663 375
rect 9701 363 9735 375
rect 9773 363 9807 375
rect 9845 363 9879 375
rect 9917 363 9951 375
rect 9989 363 10023 375
rect 10061 363 10095 375
rect 10133 363 10167 375
rect 10205 363 10239 375
rect 10277 363 10311 375
rect 10349 363 10383 375
rect 10421 363 10455 375
rect 10493 363 10527 375
rect 10565 363 10599 375
rect 10637 363 10671 375
rect 10709 363 10743 375
rect 10781 363 10815 375
rect 10853 363 10887 375
rect 10925 363 10959 375
rect 10997 363 11031 375
rect 11069 363 11103 375
rect 11141 363 11175 375
rect 11213 363 11247 375
rect 11285 363 11319 375
rect 11357 363 11391 375
rect 11429 363 11463 375
rect 11501 363 11535 375
rect 11573 363 11607 375
rect 11645 363 11679 375
rect 11717 363 11751 375
rect 11789 363 11823 375
rect 11861 363 11895 375
rect 11933 363 11967 375
rect 12005 363 12039 375
rect 12077 363 12111 375
rect 12149 363 12183 375
rect 12221 363 12255 375
rect 12293 363 12327 375
rect 12365 363 12399 375
rect 12437 363 12471 375
rect 12509 363 12543 375
rect 12581 363 12615 375
rect 12653 363 12687 375
rect 12725 363 12759 375
rect 12797 363 12831 375
rect 12869 363 12903 375
rect 12941 363 12975 375
rect 13013 363 13047 375
rect 13085 363 13119 375
rect 13157 363 13191 375
rect 13229 363 13263 375
rect 13301 363 13335 375
rect 13373 363 13407 375
rect 13445 363 13479 375
rect 13517 363 13551 375
rect 13589 363 13623 375
rect 13661 363 13695 375
rect 13733 363 13767 375
rect 13805 363 13839 375
rect 13877 363 13911 375
rect 13949 363 13983 375
rect 14021 363 14055 375
rect 14093 363 14127 375
rect 14165 363 14199 375
rect 14237 363 14271 375
rect 14309 363 14343 375
rect 14381 363 14415 375
rect 14453 363 14487 375
rect 14525 363 14559 375
rect 14597 363 14631 375
rect 14669 363 14703 375
rect 14741 363 14775 375
rect 14907 363 15051 382
rect 51 331 229 360
rect 361 341 375 363
rect 375 341 395 363
rect 434 341 448 363
rect 448 341 468 363
rect 507 341 521 363
rect 521 341 541 363
rect 580 341 594 363
rect 594 341 614 363
rect 653 341 667 363
rect 667 341 687 363
rect 726 341 740 363
rect 740 341 760 363
rect 799 341 813 363
rect 813 341 833 363
rect 872 341 886 363
rect 886 341 906 363
rect 945 341 959 363
rect 959 341 979 363
rect 1018 341 1032 363
rect 1032 341 1052 363
rect 1091 341 1105 363
rect 1105 341 1125 363
rect 1164 341 1178 363
rect 1178 341 1198 363
rect 1237 341 1251 363
rect 1251 341 1271 363
rect 1310 341 1324 363
rect 1324 341 1344 363
rect 1383 341 1397 363
rect 1397 341 1417 363
rect 1456 341 1470 363
rect 1470 341 1490 363
rect 1529 341 1543 363
rect 1543 341 1563 363
rect 1602 341 1616 363
rect 1616 341 1636 363
rect 1675 341 1689 363
rect 1689 341 1709 363
rect 1748 341 1762 363
rect 1762 341 1782 363
rect 1821 341 1835 363
rect 1835 341 1855 363
rect 1894 341 1908 363
rect 1908 341 1928 363
rect 1967 341 1981 363
rect 1981 341 2001 363
rect 2040 341 2054 363
rect 2054 341 2074 363
rect 2113 341 2127 363
rect 2127 341 2147 363
rect 2186 341 2200 363
rect 2200 341 2220 363
rect 2259 341 2273 363
rect 2273 341 2293 363
rect 2332 341 2346 363
rect 2346 341 2366 363
rect 2405 341 2419 363
rect 2419 341 2439 363
rect 2478 341 2492 363
rect 2492 341 2512 363
rect 2551 341 2565 363
rect 2565 341 2585 363
rect 2624 341 2638 363
rect 2638 341 2658 363
rect 2697 341 2711 363
rect 2711 341 2731 363
rect 2770 341 2784 363
rect 2784 341 2804 363
rect 2843 341 2857 363
rect 2857 341 2877 363
rect 2916 341 2930 363
rect 2930 341 2950 363
rect 2989 341 3003 363
rect 3003 341 3023 363
rect 3062 341 3076 363
rect 3076 341 3096 363
rect 3135 341 3149 363
rect 3149 341 3169 363
rect 3208 341 3222 363
rect 3222 341 3242 363
rect 3281 341 3295 363
rect 3295 341 3315 363
rect 3354 341 3368 363
rect 3368 341 3388 363
rect 3427 341 3440 363
rect 3440 341 3461 363
rect 3500 341 3512 363
rect 3512 341 3534 363
rect 3573 341 3584 363
rect 3584 341 3607 363
rect 3646 341 3656 363
rect 3656 341 3680 363
rect 3719 341 3728 363
rect 3728 341 3753 363
rect 3792 341 3800 363
rect 3800 341 3826 363
rect 3865 341 3872 363
rect 3872 341 3899 363
rect 3938 341 3944 363
rect 3944 341 3972 363
rect 4011 341 4016 363
rect 4016 341 4045 363
rect 4084 341 4088 363
rect 4088 341 4118 363
rect 4157 341 4160 363
rect 4160 341 4191 363
rect 4229 341 4232 363
rect 4232 341 4263 363
rect 4301 341 4304 363
rect 4304 341 4335 363
rect 4373 341 4376 363
rect 4376 341 4407 363
rect 4445 341 4448 363
rect 4448 341 4479 363
rect 4517 341 4520 363
rect 4520 341 4551 363
rect 4589 341 4592 363
rect 4592 341 4623 363
rect 4661 341 4664 363
rect 4664 341 4695 363
rect 4733 341 4736 363
rect 4736 341 4767 363
rect 4805 341 4808 363
rect 4808 341 4839 363
rect 4877 341 4880 363
rect 4880 341 4911 363
rect 4949 341 4952 363
rect 4952 341 4983 363
rect 5021 341 5024 363
rect 5024 341 5055 363
rect 5093 341 5096 363
rect 5096 341 5127 363
rect 5165 341 5168 363
rect 5168 341 5199 363
rect 5237 341 5240 363
rect 5240 341 5271 363
rect 5309 341 5312 363
rect 5312 341 5343 363
rect 5381 341 5384 363
rect 5384 341 5415 363
rect 5453 341 5456 363
rect 5456 341 5487 363
rect 5525 341 5528 363
rect 5528 341 5559 363
rect 5597 341 5600 363
rect 5600 341 5631 363
rect 5669 341 5672 363
rect 5672 341 5703 363
rect 5741 341 5744 363
rect 5744 341 5775 363
rect 5813 341 5816 363
rect 5816 341 5847 363
rect 5885 341 5888 363
rect 5888 341 5919 363
rect 5957 341 5960 363
rect 5960 341 5991 363
rect 6029 341 6032 363
rect 6032 341 6063 363
rect 6101 341 6104 363
rect 6104 341 6135 363
rect 6173 341 6176 363
rect 6176 341 6207 363
rect 6245 341 6248 363
rect 6248 341 6279 363
rect 6317 341 6320 363
rect 6320 341 6351 363
rect 6389 341 6392 363
rect 6392 341 6423 363
rect 6461 341 6464 363
rect 6464 341 6495 363
rect 6533 341 6536 363
rect 6536 341 6567 363
rect 6605 341 6608 363
rect 6608 341 6639 363
rect 6677 341 6680 363
rect 6680 341 6711 363
rect 6749 341 6752 363
rect 6752 341 6783 363
rect 6821 341 6824 363
rect 6824 341 6855 363
rect 6893 341 6896 363
rect 6896 341 6927 363
rect 6965 341 6968 363
rect 6968 341 6999 363
rect 7037 341 7040 363
rect 7040 341 7071 363
rect 7109 341 7112 363
rect 7112 341 7143 363
rect 7181 341 7184 363
rect 7184 341 7215 363
rect 7253 341 7256 363
rect 7256 341 7287 363
rect 7325 341 7328 363
rect 7328 341 7359 363
rect 7397 341 7400 363
rect 7400 341 7431 363
rect 7469 341 7472 363
rect 7472 341 7503 363
rect 7541 341 7544 363
rect 7544 341 7575 363
rect 7613 341 7616 363
rect 7616 341 7647 363
rect 7685 341 7688 363
rect 7688 341 7719 363
rect 7757 341 7760 363
rect 7760 341 7791 363
rect 7829 341 7832 363
rect 7832 341 7863 363
rect 7901 341 7904 363
rect 7904 341 7935 363
rect 7973 341 7976 363
rect 7976 341 8007 363
rect 8045 341 8048 363
rect 8048 341 8079 363
rect 8117 341 8120 363
rect 8120 341 8151 363
rect 8189 341 8192 363
rect 8192 341 8223 363
rect 8261 341 8264 363
rect 8264 341 8295 363
rect 8333 341 8336 363
rect 8336 341 8367 363
rect 8405 341 8408 363
rect 8408 341 8439 363
rect 8477 341 8480 363
rect 8480 341 8511 363
rect 8549 341 8552 363
rect 8552 341 8583 363
rect 8621 341 8624 363
rect 8624 341 8655 363
rect 8693 341 8696 363
rect 8696 341 8727 363
rect 8765 341 8768 363
rect 8768 341 8799 363
rect 8837 341 8840 363
rect 8840 341 8871 363
rect 8909 341 8912 363
rect 8912 341 8943 363
rect 8981 341 8984 363
rect 8984 341 9015 363
rect 9053 341 9056 363
rect 9056 341 9087 363
rect 9125 341 9128 363
rect 9128 341 9159 363
rect 9197 341 9200 363
rect 9200 341 9231 363
rect 9269 341 9272 363
rect 9272 341 9303 363
rect 9341 341 9344 363
rect 9344 341 9375 363
rect 9413 341 9416 363
rect 9416 341 9447 363
rect 9485 341 9488 363
rect 9488 341 9519 363
rect 9557 341 9560 363
rect 9560 341 9591 363
rect 9629 341 9632 363
rect 9632 341 9663 363
rect 9701 341 9704 363
rect 9704 341 9735 363
rect 9773 341 9776 363
rect 9776 341 9807 363
rect 9845 341 9848 363
rect 9848 341 9879 363
rect 9917 341 9920 363
rect 9920 341 9951 363
rect 9989 341 9992 363
rect 9992 341 10023 363
rect 10061 341 10064 363
rect 10064 341 10095 363
rect 10133 341 10136 363
rect 10136 341 10167 363
rect 10205 341 10208 363
rect 10208 341 10239 363
rect 10277 341 10280 363
rect 10280 341 10311 363
rect 10349 341 10352 363
rect 10352 341 10383 363
rect 10421 341 10424 363
rect 10424 341 10455 363
rect 10493 341 10496 363
rect 10496 341 10527 363
rect 10565 341 10568 363
rect 10568 341 10599 363
rect 10637 341 10640 363
rect 10640 341 10671 363
rect 10709 341 10712 363
rect 10712 341 10743 363
rect 10781 341 10784 363
rect 10784 341 10815 363
rect 10853 341 10856 363
rect 10856 341 10887 363
rect 10925 341 10928 363
rect 10928 341 10959 363
rect 10997 341 11000 363
rect 11000 341 11031 363
rect 11069 341 11072 363
rect 11072 341 11103 363
rect 11141 341 11144 363
rect 11144 341 11175 363
rect 11213 341 11216 363
rect 11216 341 11247 363
rect 11285 341 11288 363
rect 11288 341 11319 363
rect 11357 341 11360 363
rect 11360 341 11391 363
rect 11429 341 11432 363
rect 11432 341 11463 363
rect 11501 341 11504 363
rect 11504 341 11535 363
rect 11573 341 11576 363
rect 11576 341 11607 363
rect 11645 341 11648 363
rect 11648 341 11679 363
rect 11717 341 11720 363
rect 11720 341 11751 363
rect 11789 341 11792 363
rect 11792 341 11823 363
rect 11861 341 11864 363
rect 11864 341 11895 363
rect 11933 341 11936 363
rect 11936 341 11967 363
rect 12005 341 12008 363
rect 12008 341 12039 363
rect 12077 341 12080 363
rect 12080 341 12111 363
rect 12149 341 12152 363
rect 12152 341 12183 363
rect 12221 341 12224 363
rect 12224 341 12255 363
rect 12293 341 12296 363
rect 12296 341 12327 363
rect 12365 341 12368 363
rect 12368 341 12399 363
rect 12437 341 12440 363
rect 12440 341 12471 363
rect 12509 341 12512 363
rect 12512 341 12543 363
rect 12581 341 12584 363
rect 12584 341 12615 363
rect 12653 341 12656 363
rect 12656 341 12687 363
rect 12725 341 12728 363
rect 12728 341 12759 363
rect 12797 341 12800 363
rect 12800 341 12831 363
rect 12869 341 12872 363
rect 12872 341 12903 363
rect 12941 341 12944 363
rect 12944 341 12975 363
rect 13013 341 13016 363
rect 13016 341 13047 363
rect 13085 341 13088 363
rect 13088 341 13119 363
rect 13157 341 13160 363
rect 13160 341 13191 363
rect 13229 341 13232 363
rect 13232 341 13263 363
rect 13301 341 13304 363
rect 13304 341 13335 363
rect 13373 341 13376 363
rect 13376 341 13407 363
rect 13445 341 13448 363
rect 13448 341 13479 363
rect 13517 341 13520 363
rect 13520 341 13551 363
rect 13589 341 13592 363
rect 13592 341 13623 363
rect 13661 341 13664 363
rect 13664 341 13695 363
rect 13733 341 13736 363
rect 13736 341 13767 363
rect 13805 341 13808 363
rect 13808 341 13839 363
rect 13877 341 13880 363
rect 13880 341 13911 363
rect 13949 341 13952 363
rect 13952 341 13983 363
rect 14021 341 14024 363
rect 14024 341 14055 363
rect 14093 341 14096 363
rect 14096 341 14127 363
rect 14165 341 14168 363
rect 14168 341 14199 363
rect 14237 341 14240 363
rect 14240 341 14271 363
rect 14309 341 14312 363
rect 14312 341 14343 363
rect 14381 341 14384 363
rect 14384 341 14415 363
rect 14453 341 14456 363
rect 14456 341 14487 363
rect 14525 341 14528 363
rect 14528 341 14559 363
rect 14597 341 14600 363
rect 14600 341 14631 363
rect 14669 341 14672 363
rect 14672 341 14703 363
rect 14741 341 14744 363
rect 14744 341 14775 363
rect 14907 348 14922 363
rect 14922 348 14960 363
rect 14960 348 14994 363
rect 14994 348 15051 363
rect 15051 348 15085 382
<< metal1 >>
rect 39 5111 15097 5118
rect 39 5077 361 5111
rect 395 5077 434 5111
rect 468 5077 507 5111
rect 541 5077 580 5111
rect 614 5077 653 5111
rect 687 5077 726 5111
rect 760 5077 799 5111
rect 833 5077 872 5111
rect 906 5077 945 5111
rect 979 5077 1018 5111
rect 1052 5077 1091 5111
rect 1125 5077 1164 5111
rect 1198 5077 1237 5111
rect 1271 5077 1310 5111
rect 1344 5077 1383 5111
rect 1417 5077 1456 5111
rect 1490 5077 1529 5111
rect 1563 5077 1602 5111
rect 1636 5077 1675 5111
rect 1709 5077 1748 5111
rect 1782 5077 1821 5111
rect 1855 5077 1894 5111
rect 1928 5077 1967 5111
rect 2001 5077 2040 5111
rect 2074 5077 2113 5111
rect 2147 5077 2186 5111
rect 2220 5077 2259 5111
rect 2293 5077 2332 5111
rect 2366 5077 2405 5111
rect 2439 5077 2478 5111
rect 2512 5077 2551 5111
rect 2585 5077 2624 5111
rect 2658 5077 2697 5111
rect 2731 5077 2770 5111
rect 2804 5077 2843 5111
rect 2877 5077 2916 5111
rect 2950 5077 2989 5111
rect 3023 5077 3062 5111
rect 3096 5077 3135 5111
rect 3169 5077 3208 5111
rect 3242 5077 3281 5111
rect 3315 5077 3354 5111
rect 3388 5077 3427 5111
rect 3461 5077 3500 5111
rect 3534 5077 3573 5111
rect 3607 5077 3646 5111
rect 3680 5077 3719 5111
rect 3753 5077 3792 5111
rect 3826 5077 3865 5111
rect 3899 5077 3938 5111
rect 3972 5077 4011 5111
rect 4045 5077 4084 5111
rect 4118 5077 4157 5111
rect 4191 5077 4229 5111
rect 4263 5077 4301 5111
rect 4335 5077 4373 5111
rect 4407 5077 4445 5111
rect 4479 5077 4517 5111
rect 4551 5077 4589 5111
rect 4623 5077 4661 5111
rect 4695 5077 4733 5111
rect 4767 5077 4805 5111
rect 4839 5077 4877 5111
rect 4911 5077 4949 5111
rect 4983 5077 5021 5111
rect 5055 5077 5093 5111
rect 5127 5077 5165 5111
rect 5199 5077 5237 5111
rect 5271 5077 5309 5111
rect 5343 5077 5381 5111
rect 5415 5077 5453 5111
rect 5487 5077 5525 5111
rect 5559 5077 5597 5111
rect 5631 5077 5669 5111
rect 5703 5077 5741 5111
rect 5775 5077 5813 5111
rect 5847 5077 5885 5111
rect 5919 5077 5957 5111
rect 5991 5077 6029 5111
rect 6063 5077 6101 5111
rect 6135 5077 6173 5111
rect 6207 5077 6245 5111
rect 6279 5077 6317 5111
rect 6351 5077 6389 5111
rect 6423 5077 6461 5111
rect 6495 5077 6533 5111
rect 6567 5077 6605 5111
rect 6639 5077 6677 5111
rect 6711 5077 6749 5111
rect 6783 5077 6821 5111
rect 6855 5077 6893 5111
rect 6927 5077 6965 5111
rect 6999 5077 7037 5111
rect 7071 5077 7109 5111
rect 7143 5077 7181 5111
rect 7215 5077 7253 5111
rect 7287 5077 7325 5111
rect 7359 5077 7397 5111
rect 7431 5077 7469 5111
rect 7503 5077 7541 5111
rect 7575 5077 7613 5111
rect 7647 5077 7685 5111
rect 7719 5077 7757 5111
rect 7791 5077 7829 5111
rect 7863 5077 7901 5111
rect 7935 5077 7973 5111
rect 8007 5077 8045 5111
rect 8079 5077 8117 5111
rect 8151 5077 8189 5111
rect 8223 5077 8261 5111
rect 8295 5077 8333 5111
rect 8367 5077 8405 5111
rect 8439 5077 8477 5111
rect 8511 5077 8549 5111
rect 8583 5077 8621 5111
rect 8655 5077 8693 5111
rect 8727 5077 8765 5111
rect 8799 5077 8837 5111
rect 8871 5077 8909 5111
rect 8943 5077 8981 5111
rect 9015 5077 9053 5111
rect 9087 5077 9125 5111
rect 9159 5077 9197 5111
rect 9231 5077 9269 5111
rect 9303 5077 9341 5111
rect 9375 5077 9413 5111
rect 9447 5077 9485 5111
rect 9519 5077 9557 5111
rect 9591 5077 9629 5111
rect 9663 5077 9701 5111
rect 9735 5077 9773 5111
rect 9807 5077 9845 5111
rect 9879 5077 9917 5111
rect 9951 5077 9989 5111
rect 10023 5077 10061 5111
rect 10095 5077 10133 5111
rect 10167 5077 10205 5111
rect 10239 5077 10277 5111
rect 10311 5077 10349 5111
rect 10383 5077 10421 5111
rect 10455 5077 10493 5111
rect 10527 5077 10565 5111
rect 10599 5077 10637 5111
rect 10671 5077 10709 5111
rect 10743 5077 10781 5111
rect 10815 5077 10853 5111
rect 10887 5077 10925 5111
rect 10959 5077 10997 5111
rect 11031 5077 11069 5111
rect 11103 5077 11141 5111
rect 11175 5077 11213 5111
rect 11247 5077 11285 5111
rect 11319 5077 11357 5111
rect 11391 5077 11429 5111
rect 11463 5077 11501 5111
rect 11535 5077 11573 5111
rect 11607 5077 11645 5111
rect 11679 5077 11717 5111
rect 11751 5077 11789 5111
rect 11823 5077 11861 5111
rect 11895 5077 11933 5111
rect 11967 5077 12005 5111
rect 12039 5077 12077 5111
rect 12111 5077 12149 5111
rect 12183 5077 12221 5111
rect 12255 5077 12293 5111
rect 12327 5077 12365 5111
rect 12399 5077 12437 5111
rect 12471 5077 12509 5111
rect 12543 5077 12581 5111
rect 12615 5077 12653 5111
rect 12687 5077 12725 5111
rect 12759 5077 12797 5111
rect 12831 5077 12869 5111
rect 12903 5077 12941 5111
rect 12975 5077 13013 5111
rect 13047 5077 13085 5111
rect 13119 5077 13157 5111
rect 13191 5077 13229 5111
rect 13263 5077 13301 5111
rect 13335 5077 13373 5111
rect 13407 5077 13445 5111
rect 13479 5077 13517 5111
rect 13551 5077 13589 5111
rect 13623 5077 13661 5111
rect 13695 5077 13733 5111
rect 13767 5077 13805 5111
rect 13839 5077 13877 5111
rect 13911 5077 13949 5111
rect 13983 5077 14021 5111
rect 14055 5077 14093 5111
rect 14127 5077 14165 5111
rect 14199 5077 14237 5111
rect 14271 5077 14309 5111
rect 14343 5077 14381 5111
rect 14415 5077 14453 5111
rect 14487 5077 14525 5111
rect 14559 5077 14597 5111
rect 14631 5077 14669 5111
rect 14703 5077 14741 5111
rect 14775 5077 15097 5111
rect 39 5062 15097 5077
rect 39 5045 14907 5062
rect 39 331 51 5045
rect 229 5035 14907 5045
rect 229 5029 361 5035
rect 229 4995 269 5029
rect 303 5001 361 5029
rect 395 5001 434 5035
rect 468 5001 507 5035
rect 541 5001 580 5035
rect 614 5001 653 5035
rect 687 5001 726 5035
rect 760 5001 799 5035
rect 833 5001 872 5035
rect 906 5001 945 5035
rect 979 5001 1018 5035
rect 1052 5001 1091 5035
rect 1125 5001 1164 5035
rect 1198 5001 1237 5035
rect 1271 5001 1310 5035
rect 1344 5001 1383 5035
rect 1417 5001 1456 5035
rect 1490 5001 1529 5035
rect 1563 5001 1602 5035
rect 1636 5001 1675 5035
rect 1709 5001 1748 5035
rect 1782 5001 1821 5035
rect 1855 5001 1894 5035
rect 1928 5001 1967 5035
rect 2001 5001 2040 5035
rect 2074 5001 2113 5035
rect 2147 5001 2186 5035
rect 2220 5001 2259 5035
rect 2293 5001 2332 5035
rect 2366 5001 2405 5035
rect 2439 5001 2478 5035
rect 2512 5001 2551 5035
rect 2585 5001 2624 5035
rect 2658 5001 2697 5035
rect 2731 5001 2770 5035
rect 2804 5001 2843 5035
rect 2877 5001 2916 5035
rect 2950 5001 2989 5035
rect 3023 5001 3062 5035
rect 3096 5001 3135 5035
rect 3169 5001 3208 5035
rect 3242 5001 3281 5035
rect 3315 5001 3354 5035
rect 3388 5001 3427 5035
rect 3461 5001 3500 5035
rect 3534 5001 3573 5035
rect 3607 5001 3646 5035
rect 3680 5001 3719 5035
rect 3753 5001 3792 5035
rect 3826 5001 3865 5035
rect 3899 5001 3938 5035
rect 3972 5001 4011 5035
rect 4045 5001 4084 5035
rect 4118 5001 4157 5035
rect 4191 5001 4229 5035
rect 4263 5001 4301 5035
rect 4335 5001 4373 5035
rect 4407 5001 4445 5035
rect 4479 5001 4517 5035
rect 4551 5001 4589 5035
rect 4623 5001 4661 5035
rect 4695 5001 4733 5035
rect 4767 5001 4805 5035
rect 4839 5001 4877 5035
rect 4911 5001 4949 5035
rect 4983 5001 5021 5035
rect 5055 5001 5093 5035
rect 5127 5001 5165 5035
rect 5199 5001 5237 5035
rect 5271 5001 5309 5035
rect 5343 5001 5381 5035
rect 5415 5001 5453 5035
rect 5487 5001 5525 5035
rect 5559 5001 5597 5035
rect 5631 5001 5669 5035
rect 5703 5001 5741 5035
rect 5775 5001 5813 5035
rect 5847 5001 5885 5035
rect 5919 5001 5957 5035
rect 5991 5001 6029 5035
rect 6063 5001 6101 5035
rect 6135 5001 6173 5035
rect 6207 5001 6245 5035
rect 6279 5001 6317 5035
rect 6351 5001 6389 5035
rect 6423 5001 6461 5035
rect 6495 5001 6533 5035
rect 6567 5001 6605 5035
rect 6639 5001 6677 5035
rect 6711 5001 6749 5035
rect 6783 5001 6821 5035
rect 6855 5001 6893 5035
rect 6927 5001 6965 5035
rect 6999 5001 7037 5035
rect 7071 5001 7109 5035
rect 7143 5001 7181 5035
rect 7215 5001 7253 5035
rect 7287 5001 7325 5035
rect 7359 5001 7397 5035
rect 7431 5001 7469 5035
rect 7503 5001 7541 5035
rect 7575 5001 7613 5035
rect 7647 5001 7685 5035
rect 7719 5001 7757 5035
rect 7791 5001 7829 5035
rect 7863 5001 7901 5035
rect 7935 5001 7973 5035
rect 8007 5001 8045 5035
rect 8079 5001 8117 5035
rect 8151 5001 8189 5035
rect 8223 5001 8261 5035
rect 8295 5001 8333 5035
rect 8367 5001 8405 5035
rect 8439 5001 8477 5035
rect 8511 5001 8549 5035
rect 8583 5001 8621 5035
rect 8655 5001 8693 5035
rect 8727 5001 8765 5035
rect 8799 5001 8837 5035
rect 8871 5001 8909 5035
rect 8943 5001 8981 5035
rect 9015 5001 9053 5035
rect 9087 5001 9125 5035
rect 9159 5001 9197 5035
rect 9231 5001 9269 5035
rect 9303 5001 9341 5035
rect 9375 5001 9413 5035
rect 9447 5001 9485 5035
rect 9519 5001 9557 5035
rect 9591 5001 9629 5035
rect 9663 5001 9701 5035
rect 9735 5001 9773 5035
rect 9807 5001 9845 5035
rect 9879 5001 9917 5035
rect 9951 5001 9989 5035
rect 10023 5001 10061 5035
rect 10095 5001 10133 5035
rect 10167 5001 10205 5035
rect 10239 5001 10277 5035
rect 10311 5001 10349 5035
rect 10383 5001 10421 5035
rect 10455 5001 10493 5035
rect 10527 5001 10565 5035
rect 10599 5001 10637 5035
rect 10671 5001 10709 5035
rect 10743 5001 10781 5035
rect 10815 5001 10853 5035
rect 10887 5001 10925 5035
rect 10959 5001 10997 5035
rect 11031 5001 11069 5035
rect 11103 5001 11141 5035
rect 11175 5001 11213 5035
rect 11247 5001 11285 5035
rect 11319 5001 11357 5035
rect 11391 5001 11429 5035
rect 11463 5001 11501 5035
rect 11535 5001 11573 5035
rect 11607 5001 11645 5035
rect 11679 5001 11717 5035
rect 11751 5001 11789 5035
rect 11823 5001 11861 5035
rect 11895 5001 11933 5035
rect 11967 5001 12005 5035
rect 12039 5001 12077 5035
rect 12111 5001 12149 5035
rect 12183 5001 12221 5035
rect 12255 5001 12293 5035
rect 12327 5001 12365 5035
rect 12399 5001 12437 5035
rect 12471 5001 12509 5035
rect 12543 5001 12581 5035
rect 12615 5001 12653 5035
rect 12687 5001 12725 5035
rect 12759 5001 12797 5035
rect 12831 5001 12869 5035
rect 12903 5001 12941 5035
rect 12975 5001 13013 5035
rect 13047 5001 13085 5035
rect 13119 5001 13157 5035
rect 13191 5001 13229 5035
rect 13263 5001 13301 5035
rect 13335 5001 13373 5035
rect 13407 5001 13445 5035
rect 13479 5001 13517 5035
rect 13551 5001 13589 5035
rect 13623 5001 13661 5035
rect 13695 5001 13733 5035
rect 13767 5001 13805 5035
rect 13839 5001 13877 5035
rect 13911 5001 13949 5035
rect 13983 5001 14021 5035
rect 14055 5001 14093 5035
rect 14127 5001 14165 5035
rect 14199 5001 14237 5035
rect 14271 5001 14309 5035
rect 14343 5001 14381 5035
rect 14415 5001 14453 5035
rect 14487 5001 14525 5035
rect 14559 5001 14597 5035
rect 14631 5001 14669 5035
rect 14703 5001 14741 5035
rect 14775 5030 14907 5035
rect 14775 5001 14832 5030
rect 303 4996 14832 5001
rect 14866 4996 14907 5030
rect 303 4995 14907 4996
rect 229 4959 14907 4995
rect 229 4956 361 4959
rect 229 4922 269 4956
rect 303 4925 361 4956
rect 395 4925 434 4959
rect 468 4925 507 4959
rect 541 4925 580 4959
rect 614 4925 653 4959
rect 687 4925 726 4959
rect 760 4925 799 4959
rect 833 4925 872 4959
rect 906 4925 945 4959
rect 979 4925 1018 4959
rect 1052 4925 1091 4959
rect 1125 4925 1164 4959
rect 1198 4925 1237 4959
rect 1271 4925 1310 4959
rect 1344 4925 1383 4959
rect 1417 4925 1456 4959
rect 1490 4925 1529 4959
rect 1563 4925 1602 4959
rect 1636 4925 1675 4959
rect 1709 4925 1748 4959
rect 1782 4925 1821 4959
rect 1855 4925 1894 4959
rect 1928 4925 1967 4959
rect 2001 4925 2040 4959
rect 2074 4925 2113 4959
rect 2147 4925 2186 4959
rect 2220 4925 2259 4959
rect 2293 4925 2332 4959
rect 2366 4925 2405 4959
rect 2439 4925 2478 4959
rect 2512 4925 2551 4959
rect 2585 4925 2624 4959
rect 2658 4925 2697 4959
rect 2731 4925 2770 4959
rect 2804 4925 2843 4959
rect 2877 4925 2916 4959
rect 2950 4925 2989 4959
rect 3023 4925 3062 4959
rect 3096 4925 3135 4959
rect 3169 4925 3208 4959
rect 3242 4925 3281 4959
rect 3315 4925 3354 4959
rect 3388 4925 3427 4959
rect 3461 4925 3500 4959
rect 3534 4925 3573 4959
rect 3607 4925 3646 4959
rect 3680 4925 3719 4959
rect 3753 4925 3792 4959
rect 3826 4925 3865 4959
rect 3899 4925 3938 4959
rect 3972 4925 4011 4959
rect 4045 4925 4084 4959
rect 4118 4925 4157 4959
rect 4191 4925 4229 4959
rect 4263 4925 4301 4959
rect 4335 4925 4373 4959
rect 4407 4925 4445 4959
rect 4479 4925 4517 4959
rect 4551 4925 4589 4959
rect 4623 4925 4661 4959
rect 4695 4925 4733 4959
rect 4767 4925 4805 4959
rect 4839 4925 4877 4959
rect 4911 4925 4949 4959
rect 4983 4925 5021 4959
rect 5055 4925 5093 4959
rect 5127 4925 5165 4959
rect 5199 4925 5237 4959
rect 5271 4925 5309 4959
rect 5343 4925 5381 4959
rect 5415 4925 5453 4959
rect 5487 4925 5525 4959
rect 5559 4925 5597 4959
rect 5631 4925 5669 4959
rect 5703 4925 5741 4959
rect 5775 4925 5813 4959
rect 5847 4925 5885 4959
rect 5919 4925 5957 4959
rect 5991 4925 6029 4959
rect 6063 4925 6101 4959
rect 6135 4925 6173 4959
rect 6207 4925 6245 4959
rect 6279 4925 6317 4959
rect 6351 4925 6389 4959
rect 6423 4925 6461 4959
rect 6495 4925 6533 4959
rect 6567 4925 6605 4959
rect 6639 4925 6677 4959
rect 6711 4925 6749 4959
rect 6783 4925 6821 4959
rect 6855 4925 6893 4959
rect 6927 4925 6965 4959
rect 6999 4925 7037 4959
rect 7071 4925 7109 4959
rect 7143 4925 7181 4959
rect 7215 4925 7253 4959
rect 7287 4925 7325 4959
rect 7359 4925 7397 4959
rect 7431 4925 7469 4959
rect 7503 4925 7541 4959
rect 7575 4925 7613 4959
rect 7647 4925 7685 4959
rect 7719 4925 7757 4959
rect 7791 4925 7829 4959
rect 7863 4925 7901 4959
rect 7935 4925 7973 4959
rect 8007 4925 8045 4959
rect 8079 4925 8117 4959
rect 8151 4925 8189 4959
rect 8223 4925 8261 4959
rect 8295 4925 8333 4959
rect 8367 4925 8405 4959
rect 8439 4925 8477 4959
rect 8511 4925 8549 4959
rect 8583 4925 8621 4959
rect 8655 4925 8693 4959
rect 8727 4925 8765 4959
rect 8799 4925 8837 4959
rect 8871 4925 8909 4959
rect 8943 4925 8981 4959
rect 9015 4925 9053 4959
rect 9087 4925 9125 4959
rect 9159 4925 9197 4959
rect 9231 4925 9269 4959
rect 9303 4925 9341 4959
rect 9375 4925 9413 4959
rect 9447 4925 9485 4959
rect 9519 4925 9557 4959
rect 9591 4925 9629 4959
rect 9663 4925 9701 4959
rect 9735 4925 9773 4959
rect 9807 4925 9845 4959
rect 9879 4925 9917 4959
rect 9951 4925 9989 4959
rect 10023 4925 10061 4959
rect 10095 4925 10133 4959
rect 10167 4925 10205 4959
rect 10239 4925 10277 4959
rect 10311 4925 10349 4959
rect 10383 4925 10421 4959
rect 10455 4925 10493 4959
rect 10527 4925 10565 4959
rect 10599 4925 10637 4959
rect 10671 4925 10709 4959
rect 10743 4925 10781 4959
rect 10815 4925 10853 4959
rect 10887 4925 10925 4959
rect 10959 4925 10997 4959
rect 11031 4925 11069 4959
rect 11103 4925 11141 4959
rect 11175 4925 11213 4959
rect 11247 4925 11285 4959
rect 11319 4925 11357 4959
rect 11391 4925 11429 4959
rect 11463 4925 11501 4959
rect 11535 4925 11573 4959
rect 11607 4925 11645 4959
rect 11679 4925 11717 4959
rect 11751 4925 11789 4959
rect 11823 4925 11861 4959
rect 11895 4925 11933 4959
rect 11967 4925 12005 4959
rect 12039 4925 12077 4959
rect 12111 4925 12149 4959
rect 12183 4925 12221 4959
rect 12255 4925 12293 4959
rect 12327 4925 12365 4959
rect 12399 4925 12437 4959
rect 12471 4925 12509 4959
rect 12543 4925 12581 4959
rect 12615 4925 12653 4959
rect 12687 4925 12725 4959
rect 12759 4925 12797 4959
rect 12831 4925 12869 4959
rect 12903 4925 12941 4959
rect 12975 4925 13013 4959
rect 13047 4925 13085 4959
rect 13119 4925 13157 4959
rect 13191 4925 13229 4959
rect 13263 4925 13301 4959
rect 13335 4925 13373 4959
rect 13407 4925 13445 4959
rect 13479 4925 13517 4959
rect 13551 4925 13589 4959
rect 13623 4925 13661 4959
rect 13695 4925 13733 4959
rect 13767 4925 13805 4959
rect 13839 4925 13877 4959
rect 13911 4925 13949 4959
rect 13983 4925 14021 4959
rect 14055 4925 14093 4959
rect 14127 4925 14165 4959
rect 14199 4925 14237 4959
rect 14271 4925 14309 4959
rect 14343 4925 14381 4959
rect 14415 4925 14453 4959
rect 14487 4925 14525 4959
rect 14559 4925 14597 4959
rect 14631 4925 14669 4959
rect 14703 4925 14741 4959
rect 14775 4958 14907 4959
rect 14775 4925 14832 4958
rect 303 4924 14832 4925
rect 14866 4924 14907 4958
rect 303 4922 14907 4924
rect 229 4918 14907 4922
rect 229 4886 759 4918
tri 759 4886 791 4918 nw
tri 14335 4886 14367 4918 ne
rect 14367 4886 14907 4918
rect 229 4883 725 4886
rect 229 4849 269 4883
rect 303 4852 725 4883
tri 725 4852 759 4886 nw
tri 14367 4852 14401 4886 ne
rect 14401 4852 14832 4886
rect 14866 4852 14907 4886
rect 303 4849 687 4852
rect 229 4814 687 4849
tri 687 4814 725 4852 nw
tri 14401 4814 14439 4852 ne
rect 14439 4814 14907 4852
rect 229 4810 653 4814
rect 229 4776 269 4810
rect 303 4780 653 4810
tri 653 4780 687 4814 nw
tri 14439 4780 14473 4814 ne
rect 14473 4780 14832 4814
rect 14866 4780 14907 4814
rect 303 4776 615 4780
rect 229 4742 615 4776
tri 615 4742 653 4780 nw
tri 14473 4742 14511 4780 ne
rect 14511 4742 14907 4780
rect 229 4737 581 4742
rect 229 4703 269 4737
rect 303 4708 581 4737
tri 581 4708 615 4742 nw
tri 14511 4708 14545 4742 ne
rect 14545 4708 14832 4742
rect 14866 4708 14907 4742
rect 303 4703 543 4708
rect 229 4670 543 4703
tri 543 4670 581 4708 nw
tri 14545 4670 14583 4708 ne
rect 14583 4670 14907 4708
rect 229 4664 509 4670
rect 229 4630 269 4664
rect 303 4636 509 4664
tri 509 4636 543 4670 nw
tri 14583 4636 14617 4670 ne
rect 14617 4636 14832 4670
rect 14866 4636 14907 4670
rect 303 4630 491 4636
rect 229 4618 491 4630
tri 491 4618 509 4636 nw
tri 14617 4618 14635 4636 ne
rect 14635 4618 14907 4636
rect 229 4606 479 4618
tri 479 4606 491 4618 nw
tri 621 4606 633 4618 se
rect 633 4606 14502 4618
rect 229 4591 373 4606
rect 229 4557 269 4591
rect 303 4557 373 4591
rect 229 4518 373 4557
rect 229 4484 269 4518
rect 303 4500 373 4518
tri 373 4500 479 4606 nw
tri 517 4502 621 4606 se
rect 621 4502 709 4606
rect 517 4500 709 4502
rect 14207 4572 14246 4606
rect 14280 4572 14319 4606
rect 14353 4572 14392 4606
rect 14426 4598 14502 4606
tri 14502 4598 14522 4618 sw
tri 14635 4598 14655 4618 ne
rect 14655 4598 14907 4618
rect 14426 4572 14522 4598
rect 14207 4564 14522 4572
tri 14522 4564 14556 4598 sw
tri 14655 4564 14689 4598 ne
rect 14689 4564 14832 4598
rect 14866 4564 14907 4598
rect 14207 4534 14556 4564
rect 14207 4500 14246 4534
rect 14280 4500 14319 4534
rect 14353 4500 14392 4534
rect 14426 4526 14556 4534
tri 14556 4526 14594 4564 sw
tri 14689 4526 14727 4564 ne
rect 14727 4526 14907 4564
rect 14426 4502 14594 4526
tri 14594 4502 14618 4526 sw
rect 14426 4500 14618 4502
rect 303 4492 365 4500
tri 365 4492 373 4500 nw
rect 303 4484 329 4492
rect 229 4445 329 4484
tri 329 4456 365 4492 nw
rect 517 4488 14618 4500
tri 14727 4492 14761 4526 ne
rect 14761 4492 14832 4526
rect 14866 4492 14907 4526
rect 517 4456 946 4488
tri 946 4456 978 4488 nw
tri 14157 4468 14177 4488 ne
rect 14177 4468 14618 4488
tri 14177 4456 14189 4468 ne
rect 14189 4456 14618 4468
rect 229 4411 269 4445
rect 303 4411 329 4445
rect 229 4372 329 4411
rect 229 4338 269 4372
rect 303 4338 329 4372
rect 229 4299 329 4338
rect 229 4265 269 4299
rect 303 4265 329 4299
rect 229 4226 329 4265
rect 229 4192 269 4226
rect 303 4192 329 4226
rect 229 4153 329 4192
rect 229 4119 269 4153
rect 303 4119 329 4153
rect 229 4080 329 4119
rect 229 4046 269 4080
rect 303 4046 329 4080
rect 229 4007 329 4046
rect 229 3973 269 4007
rect 303 3973 329 4007
rect 229 3934 329 3973
rect 229 3900 269 3934
rect 303 3900 329 3934
rect 229 3861 329 3900
rect 229 3827 269 3861
rect 303 3827 329 3861
rect 229 3788 329 3827
rect 229 3754 269 3788
rect 303 3754 329 3788
rect 229 3715 329 3754
rect 229 3681 269 3715
rect 303 3681 329 3715
rect 229 3642 329 3681
rect 229 3608 269 3642
rect 303 3608 329 3642
rect 229 3569 329 3608
rect 229 3535 269 3569
rect 303 3535 329 3569
rect 229 3496 329 3535
rect 229 3462 269 3496
rect 303 3462 329 3496
rect 229 3423 329 3462
rect 229 3389 269 3423
rect 303 3389 329 3423
rect 229 3350 329 3389
rect 229 3316 269 3350
rect 303 3316 329 3350
rect 229 3277 329 3316
rect 229 3243 269 3277
rect 303 3243 329 3277
rect 229 3204 329 3243
rect 229 3170 269 3204
rect 303 3170 329 3204
rect 229 3131 329 3170
rect 229 3097 269 3131
rect 303 3097 329 3131
rect 229 3058 329 3097
rect 229 3024 269 3058
rect 303 3024 329 3058
rect 229 2985 329 3024
rect 229 2951 269 2985
rect 303 2951 329 2985
rect 229 2912 329 2951
rect 229 2878 269 2912
rect 303 2878 329 2912
rect 229 2839 329 2878
rect 229 2805 269 2839
rect 303 2805 329 2839
rect 229 2766 329 2805
rect 229 2732 269 2766
rect 303 2732 329 2766
rect 229 2693 329 2732
rect 229 2659 269 2693
rect 303 2659 329 2693
rect 229 2620 329 2659
rect 229 2586 269 2620
rect 303 2586 329 2620
rect 229 2547 329 2586
rect 229 2513 269 2547
rect 303 2513 329 2547
rect 229 2474 329 2513
rect 229 2440 269 2474
rect 303 2440 329 2474
rect 229 2401 329 2440
rect 229 2367 269 2401
rect 303 2367 329 2401
rect 229 2328 329 2367
rect 229 2294 269 2328
rect 303 2294 329 2328
rect 229 2255 329 2294
rect 229 2221 269 2255
rect 303 2221 329 2255
rect 229 2182 329 2221
rect 229 2148 269 2182
rect 303 2148 329 2182
rect 229 2109 329 2148
rect 229 2075 269 2109
rect 303 2075 329 2109
rect 229 2036 329 2075
rect 229 2002 269 2036
rect 303 2002 329 2036
rect 229 1963 329 2002
rect 229 1929 269 1963
rect 303 1929 329 1963
rect 229 1890 329 1929
rect 229 1856 269 1890
rect 303 1856 329 1890
rect 229 1817 329 1856
rect 229 1783 269 1817
rect 303 1783 329 1817
rect 229 1744 329 1783
rect 229 1710 269 1744
rect 303 1710 329 1744
rect 229 1671 329 1710
rect 229 1637 269 1671
rect 303 1637 329 1671
rect 229 1598 329 1637
rect 229 1564 269 1598
rect 303 1564 329 1598
rect 229 1525 329 1564
rect 229 1491 269 1525
rect 303 1491 329 1525
rect 229 1452 329 1491
rect 229 1418 269 1452
rect 303 1418 329 1452
rect 229 1379 329 1418
rect 229 1345 269 1379
rect 303 1345 329 1379
rect 229 1306 329 1345
rect 229 1272 269 1306
rect 303 1272 329 1306
rect 229 1233 329 1272
rect 229 1199 269 1233
rect 303 1199 329 1233
rect 229 1159 329 1199
rect 229 1125 269 1159
rect 303 1125 329 1159
rect 229 1085 329 1125
rect 229 1051 269 1085
rect 303 1051 329 1085
rect 229 1011 329 1051
rect 229 977 269 1011
rect 303 977 329 1011
rect 229 937 329 977
rect 229 903 269 937
rect 303 903 329 937
rect 229 863 329 903
rect 517 4426 674 4456
rect 708 4448 938 4456
tri 938 4448 946 4456 nw
tri 14189 4448 14197 4456 ne
rect 14197 4448 14428 4456
rect 708 4445 922 4448
rect 517 4392 529 4426
rect 563 4392 601 4426
rect 635 4392 674 4426
rect 517 4351 674 4392
rect 517 4317 529 4351
rect 563 4317 601 4351
rect 635 4317 674 4351
rect 517 4276 674 4317
rect 517 4242 529 4276
rect 563 4242 601 4276
rect 635 4242 674 4276
rect 517 4201 674 4242
rect 517 4167 529 4201
rect 563 4167 601 4201
rect 635 4167 674 4201
rect 517 4126 674 4167
rect 517 4092 529 4126
rect 563 4092 601 4126
rect 635 4092 674 4126
rect 517 4052 674 4092
rect 517 4018 529 4052
rect 563 4018 601 4052
rect 635 4018 674 4052
rect 517 3978 674 4018
rect 517 3944 529 3978
rect 563 3944 601 3978
rect 635 3944 674 3978
rect 517 3904 674 3944
rect 517 3870 529 3904
rect 563 3870 601 3904
rect 635 3870 674 3904
rect 517 3794 674 3870
rect 517 3760 529 3794
rect 563 3760 601 3794
rect 635 3760 674 3794
rect 517 3720 674 3760
rect 517 3686 529 3720
rect 563 3686 601 3720
rect 635 3686 674 3720
rect 517 3646 674 3686
rect 517 3612 529 3646
rect 563 3612 601 3646
rect 635 3612 674 3646
rect 517 3572 674 3612
rect 517 3538 529 3572
rect 563 3538 601 3572
rect 635 3538 674 3572
rect 517 3498 674 3538
rect 517 3464 529 3498
rect 563 3464 601 3498
rect 635 3464 674 3498
rect 517 3424 674 3464
rect 517 3390 529 3424
rect 563 3390 601 3424
rect 635 3390 674 3424
rect 517 3350 674 3390
rect 517 3316 529 3350
rect 563 3316 601 3350
rect 635 3316 674 3350
rect 517 3276 674 3316
rect 517 3242 529 3276
rect 563 3242 601 3276
rect 635 3242 674 3276
rect 517 3202 674 3242
rect 517 3168 529 3202
rect 563 3168 601 3202
rect 635 3168 674 3202
rect 517 3128 674 3168
rect 517 3094 529 3128
rect 563 3094 601 3128
rect 635 3094 674 3128
rect 517 3054 674 3094
rect 517 3020 529 3054
rect 563 3020 601 3054
rect 635 3020 674 3054
rect 517 2980 674 3020
rect 517 2946 529 2980
rect 563 2946 601 2980
rect 635 2946 674 2980
rect 517 2906 674 2946
rect 517 2872 529 2906
rect 563 2872 601 2906
rect 635 2872 674 2906
rect 517 2832 674 2872
rect 517 2798 529 2832
rect 563 2798 601 2832
rect 635 2798 674 2832
rect 517 2758 674 2798
rect 517 2724 529 2758
rect 563 2724 601 2758
rect 635 2724 674 2758
rect 517 2684 674 2724
rect 517 2650 529 2684
rect 563 2657 601 2684
rect 635 2657 674 2684
rect 780 4432 922 4445
tri 922 4432 938 4448 nw
tri 14197 4444 14201 4448 ne
rect 14201 4444 14428 4448
tri 14201 4432 14213 4444 ne
rect 14213 4432 14428 4444
rect 780 4398 888 4432
tri 888 4398 922 4432 nw
tri 14213 4398 14247 4432 ne
rect 14247 4398 14356 4432
rect 14390 4398 14428 4432
rect 14462 4426 14618 4456
tri 14761 4454 14799 4492 ne
rect 14799 4454 14907 4492
tri 14799 4446 14807 4454 ne
rect 780 4359 849 4398
tri 849 4359 888 4398 nw
tri 14247 4359 14286 4398 ne
rect 14286 4359 14428 4398
rect 780 4325 815 4359
tri 815 4325 849 4359 nw
tri 14286 4325 14320 4359 ne
rect 14320 4325 14356 4359
rect 14390 4325 14428 4359
rect 780 2657 786 4325
tri 786 4296 815 4325 nw
tri 14320 4296 14349 4325 ne
rect 14349 4296 14428 4325
tri 14349 4295 14350 4296 ne
rect 14350 4286 14428 4296
rect 14350 4252 14356 4286
rect 14390 4252 14428 4286
rect 14350 4213 14428 4252
rect 14350 4179 14356 4213
rect 14390 4179 14428 4213
rect 14350 4140 14428 4179
rect 635 2650 646 2657
rect 517 2610 558 2650
rect 610 2610 646 2650
rect 517 2576 529 2610
rect 635 2605 646 2610
rect 563 2592 601 2605
rect 635 2592 674 2605
rect 780 2592 786 2605
rect 635 2576 646 2592
rect 517 2540 558 2576
rect 610 2540 646 2576
rect 517 2536 674 2540
rect 517 2502 529 2536
rect 563 2527 601 2536
rect 635 2527 674 2536
rect 780 2527 786 2540
rect 635 2502 646 2527
rect 517 2475 558 2502
rect 610 2475 646 2502
rect 517 2462 674 2475
rect 780 2462 786 2475
rect 517 2428 529 2462
rect 635 2428 646 2462
rect 517 2410 558 2428
rect 610 2410 646 2428
rect 517 2397 674 2410
rect 780 2397 786 2410
rect 517 2389 558 2397
rect 610 2389 646 2397
rect 517 2355 529 2389
rect 635 2355 646 2389
rect 517 2345 558 2355
rect 610 2345 646 2355
rect 517 2332 674 2345
rect 780 2332 786 2345
rect 517 2316 558 2332
rect 610 2316 646 2332
rect 517 2282 529 2316
rect 635 2282 646 2316
rect 517 2280 558 2282
rect 610 2280 646 2282
rect 517 2267 674 2280
rect 780 2267 786 2280
rect 517 2243 558 2267
rect 610 2243 646 2267
rect 517 2209 529 2243
rect 635 2215 646 2243
rect 563 2209 601 2215
rect 635 2209 674 2215
rect 517 2202 674 2209
rect 780 2202 786 2215
rect 517 2170 558 2202
rect 610 2170 646 2202
rect 517 2136 529 2170
rect 635 2150 646 2170
rect 563 2137 601 2150
rect 635 2137 674 2150
rect 780 2137 786 2150
rect 635 2136 646 2137
rect 517 2097 558 2136
rect 610 2097 646 2136
rect 517 2063 529 2097
rect 635 2085 646 2097
rect 563 2072 601 2085
rect 635 2072 674 2085
rect 780 2072 786 2085
rect 635 2063 646 2072
rect 517 2024 558 2063
rect 610 2024 646 2063
rect 517 1990 529 2024
rect 635 2020 646 2024
rect 563 2007 601 2020
rect 635 2007 674 2020
rect 780 2007 786 2020
rect 635 1990 646 2007
rect 517 1955 558 1990
rect 610 1955 646 1990
rect 517 1951 674 1955
rect 517 1917 529 1951
rect 563 1942 601 1951
rect 635 1942 674 1951
rect 780 1942 786 1955
rect 635 1917 646 1942
rect 517 1890 558 1917
rect 610 1890 646 1917
rect 517 1878 674 1890
rect 517 1844 529 1878
rect 563 1877 601 1878
rect 635 1877 674 1878
rect 780 1877 786 1890
rect 635 1844 646 1877
rect 517 1825 558 1844
rect 610 1825 646 1844
rect 517 1812 674 1825
rect 780 1812 786 1825
rect 517 1805 558 1812
rect 610 1805 646 1812
rect 517 1771 529 1805
rect 635 1771 646 1805
rect 517 1760 558 1771
rect 610 1760 646 1771
rect 517 1748 674 1760
rect 780 1748 786 1760
rect 517 1732 558 1748
rect 610 1732 646 1748
rect 517 1698 529 1732
rect 635 1698 646 1732
rect 517 1696 558 1698
rect 610 1696 646 1698
rect 517 1684 674 1696
rect 780 1684 786 1696
rect 517 1659 558 1684
rect 610 1659 646 1684
rect 517 1625 529 1659
rect 635 1632 646 1659
rect 563 1625 601 1632
rect 635 1625 674 1632
rect 517 1620 674 1625
rect 780 1620 786 1632
rect 517 1586 558 1620
rect 610 1586 646 1620
rect 517 1552 529 1586
rect 635 1568 646 1586
rect 563 1552 601 1568
rect 635 1552 674 1568
rect 517 1513 674 1552
rect 517 1479 529 1513
rect 563 1479 601 1513
rect 635 1479 674 1513
rect 517 1440 674 1479
rect 517 1406 529 1440
rect 563 1406 601 1440
rect 635 1406 674 1440
rect 517 1367 674 1406
rect 517 1333 529 1367
rect 563 1333 601 1367
rect 635 1333 674 1367
rect 517 1294 674 1333
rect 517 1260 529 1294
rect 563 1260 601 1294
rect 635 1260 674 1294
rect 517 1221 674 1260
rect 517 1187 529 1221
rect 563 1187 601 1221
rect 635 1187 674 1221
rect 517 1148 674 1187
rect 517 1114 529 1148
rect 563 1114 601 1148
rect 635 1114 674 1148
rect 517 1075 674 1114
rect 517 1041 529 1075
rect 563 1041 601 1075
rect 635 1041 674 1075
rect 517 1002 674 1041
rect 517 968 529 1002
rect 563 968 601 1002
rect 635 968 674 1002
rect 517 929 674 968
rect 517 895 529 929
rect 563 895 601 929
rect 635 895 674 929
rect 517 894 674 895
rect 780 1001 786 1568
rect 1060 4119 1252 4125
rect 1060 4067 1066 4119
rect 1118 4067 1130 4119
rect 1182 4067 1194 4119
rect 1246 4067 1252 4119
rect 1060 4064 1067 4067
rect 1101 4064 1139 4067
rect 1173 4064 1211 4067
rect 1245 4064 1252 4067
rect 1060 4054 1252 4064
rect 1060 4002 1066 4054
rect 1118 4002 1130 4054
rect 1182 4002 1194 4054
rect 1246 4002 1252 4054
rect 1060 3991 1067 4002
rect 1101 3991 1139 4002
rect 1173 3991 1211 4002
rect 1245 3991 1252 4002
rect 1060 3989 1252 3991
rect 1060 3937 1066 3989
rect 1118 3937 1130 3989
rect 1182 3937 1194 3989
rect 1246 3937 1252 3989
rect 1060 3924 1067 3937
rect 1101 3924 1139 3937
rect 1173 3924 1211 3937
rect 1245 3924 1252 3937
rect 1060 3872 1066 3924
rect 1118 3872 1130 3924
rect 1182 3872 1194 3924
rect 1246 3872 1252 3924
rect 1060 3859 1067 3872
rect 1101 3859 1139 3872
rect 1173 3859 1211 3872
rect 1245 3859 1252 3872
rect 1060 3807 1066 3859
rect 1118 3807 1130 3859
rect 1182 3807 1194 3859
rect 1246 3807 1252 3859
rect 1060 3806 1252 3807
rect 1060 3794 1067 3806
rect 1101 3794 1139 3806
rect 1173 3794 1211 3806
rect 1245 3794 1252 3806
rect 1060 3742 1066 3794
rect 1118 3742 1130 3794
rect 1182 3742 1194 3794
rect 1246 3742 1252 3794
rect 1060 3733 1252 3742
rect 1060 3729 1067 3733
rect 1101 3729 1139 3733
rect 1173 3729 1211 3733
rect 1245 3729 1252 3733
rect 1060 3677 1066 3729
rect 1118 3677 1130 3729
rect 1182 3677 1194 3729
rect 1246 3677 1252 3729
rect 1060 3664 1252 3677
rect 1060 2972 1066 3664
rect 1246 2972 1252 3664
rect 1060 2969 1067 2972
rect 1101 2969 1139 2972
rect 1173 2969 1211 2972
rect 1245 2969 1252 2972
rect 1060 2930 1252 2969
rect 1060 2896 1067 2930
rect 1101 2896 1139 2930
rect 1173 2896 1211 2930
rect 1245 2896 1252 2930
rect 1060 2857 1252 2896
rect 1060 2823 1067 2857
rect 1101 2823 1139 2857
rect 1173 2823 1211 2857
rect 1245 2823 1252 2857
rect 1060 2784 1252 2823
rect 1060 2750 1067 2784
rect 1101 2750 1139 2784
rect 1173 2750 1211 2784
rect 1245 2750 1252 2784
rect 1060 2711 1252 2750
rect 1060 2677 1067 2711
rect 1101 2677 1139 2711
rect 1173 2677 1211 2711
rect 1245 2677 1252 2711
rect 1060 2638 1252 2677
rect 1060 2604 1067 2638
rect 1101 2604 1139 2638
rect 1173 2604 1211 2638
rect 1245 2604 1252 2638
rect 1060 2565 1252 2604
rect 1060 2531 1067 2565
rect 1101 2531 1139 2565
rect 1173 2531 1211 2565
rect 1245 2531 1252 2565
rect 1060 2492 1252 2531
rect 1060 2458 1067 2492
rect 1101 2458 1139 2492
rect 1173 2458 1211 2492
rect 1245 2458 1252 2492
rect 1060 2419 1252 2458
rect 1060 2385 1067 2419
rect 1101 2385 1139 2419
rect 1173 2385 1211 2419
rect 1245 2385 1252 2419
rect 1060 2346 1252 2385
rect 1060 2312 1067 2346
rect 1101 2312 1139 2346
rect 1173 2312 1211 2346
rect 1245 2312 1252 2346
rect 1060 2273 1252 2312
rect 1060 2239 1067 2273
rect 1101 2239 1139 2273
rect 1173 2239 1211 2273
rect 1245 2239 1252 2273
rect 1060 2200 1252 2239
rect 1060 2166 1067 2200
rect 1101 2166 1139 2200
rect 1173 2166 1211 2200
rect 1245 2166 1252 2200
rect 1060 2126 1252 2166
rect 1060 2092 1067 2126
rect 1101 2092 1139 2126
rect 1173 2092 1211 2126
rect 1245 2092 1252 2126
rect 1060 2052 1252 2092
rect 1060 2018 1067 2052
rect 1101 2018 1139 2052
rect 1173 2018 1211 2052
rect 1245 2018 1252 2052
rect 1060 1978 1252 2018
rect 1060 1944 1067 1978
rect 1101 1944 1139 1978
rect 1173 1944 1211 1978
rect 1245 1944 1252 1978
rect 1060 1904 1252 1944
rect 1060 1870 1067 1904
rect 1101 1870 1139 1904
rect 1173 1870 1211 1904
rect 1245 1870 1252 1904
rect 1060 1830 1252 1870
rect 1060 1796 1067 1830
rect 1101 1796 1139 1830
rect 1173 1796 1211 1830
rect 1245 1796 1252 1830
rect 1060 1756 1252 1796
rect 1060 1722 1067 1756
rect 1101 1722 1139 1756
rect 1173 1722 1211 1756
rect 1245 1722 1252 1756
rect 1060 1682 1252 1722
rect 1060 1648 1067 1682
rect 1101 1648 1139 1682
rect 1173 1648 1211 1682
rect 1245 1648 1252 1682
rect 1060 1608 1252 1648
rect 1060 1574 1067 1608
rect 1101 1574 1139 1608
rect 1173 1574 1211 1608
rect 1245 1574 1252 1608
rect 1060 1562 1252 1574
rect 1556 4118 1748 4130
rect 1556 4092 1635 4118
rect 1669 4092 1748 4118
rect 1556 3194 1563 4092
rect 1741 3194 1748 4092
rect 1556 3182 1748 3194
rect 1556 3148 1635 3182
rect 1669 3148 1748 3182
rect 1556 3108 1748 3148
rect 1556 3074 1563 3108
rect 1597 3074 1635 3108
rect 1669 3074 1707 3108
rect 1741 3074 1748 3108
rect 1556 3028 1748 3074
rect 1556 2994 1563 3028
rect 1597 2994 1635 3028
rect 1669 2994 1707 3028
rect 1741 2994 1748 3028
rect 1556 2948 1748 2994
rect 1556 2914 1563 2948
rect 1597 2914 1635 2948
rect 1669 2914 1707 2948
rect 1741 2914 1748 2948
rect 1556 2868 1748 2914
rect 1556 2834 1563 2868
rect 1597 2834 1635 2868
rect 1669 2834 1707 2868
rect 1741 2834 1748 2868
rect 1556 2788 1748 2834
rect 1556 2754 1563 2788
rect 1597 2754 1635 2788
rect 1669 2754 1707 2788
rect 1741 2754 1748 2788
rect 1556 2708 1748 2754
rect 1556 2674 1563 2708
rect 1597 2674 1635 2708
rect 1669 2674 1707 2708
rect 1741 2674 1748 2708
rect 1556 2657 1748 2674
rect 1556 2605 1562 2657
rect 1614 2605 1626 2657
rect 1678 2605 1690 2657
rect 1742 2605 1748 2657
rect 1556 2594 1563 2605
rect 1597 2594 1635 2605
rect 1669 2594 1707 2605
rect 1741 2594 1748 2605
rect 1556 2592 1748 2594
rect 1556 2540 1562 2592
rect 1614 2540 1626 2592
rect 1678 2540 1690 2592
rect 1742 2540 1748 2592
rect 1556 2527 1635 2540
rect 1669 2527 1748 2540
rect 1556 2475 1562 2527
rect 1614 2518 1626 2527
rect 1678 2518 1690 2527
rect 1742 2475 1748 2527
rect 1556 2462 1563 2475
rect 1741 2462 1748 2475
rect 1556 2410 1562 2462
rect 1742 2410 1748 2462
rect 1556 2397 1563 2410
rect 1741 2397 1748 2410
rect 1556 2345 1562 2397
rect 1742 2345 1748 2397
rect 1556 2332 1563 2345
rect 1741 2332 1748 2345
rect 1556 2280 1562 2332
rect 1742 2280 1748 2332
rect 1556 2267 1563 2280
rect 1741 2267 1748 2280
rect 1556 2215 1562 2267
rect 1742 2215 1748 2267
rect 1556 2202 1563 2215
rect 1741 2202 1748 2215
rect 1556 2150 1562 2202
rect 1742 2150 1748 2202
rect 1556 2137 1563 2150
rect 1741 2137 1748 2150
rect 1556 2085 1562 2137
rect 1742 2085 1748 2137
rect 1556 2072 1563 2085
rect 1741 2072 1748 2085
rect 1556 2020 1562 2072
rect 1742 2020 1748 2072
rect 1556 2007 1563 2020
rect 1741 2007 1748 2020
rect 1556 1955 1562 2007
rect 1742 1955 1748 2007
rect 1556 1942 1563 1955
rect 1741 1942 1748 1955
rect 1556 1890 1562 1942
rect 1742 1890 1748 1942
rect 1556 1877 1563 1890
rect 1741 1877 1748 1890
rect 1556 1825 1562 1877
rect 1742 1825 1748 1877
rect 1556 1812 1563 1825
rect 1741 1812 1748 1825
rect 1556 1568 1562 1812
rect 1742 1568 1748 1812
rect 1556 1562 1748 1568
rect 2052 4119 2244 4125
rect 2052 4067 2058 4119
rect 2110 4067 2122 4119
rect 2174 4067 2186 4119
rect 2238 4067 2244 4119
rect 2052 4064 2059 4067
rect 2093 4064 2131 4067
rect 2165 4064 2203 4067
rect 2237 4064 2244 4067
rect 2052 4054 2244 4064
rect 2052 4002 2058 4054
rect 2110 4002 2122 4054
rect 2174 4002 2186 4054
rect 2238 4002 2244 4054
rect 2052 3991 2059 4002
rect 2093 3991 2131 4002
rect 2165 3991 2203 4002
rect 2237 3991 2244 4002
rect 2052 3989 2244 3991
rect 2052 3937 2058 3989
rect 2110 3937 2122 3989
rect 2174 3937 2186 3989
rect 2238 3937 2244 3989
rect 2052 3924 2059 3937
rect 2093 3924 2131 3937
rect 2165 3924 2203 3937
rect 2237 3924 2244 3937
rect 2052 3872 2058 3924
rect 2110 3872 2122 3924
rect 2174 3872 2186 3924
rect 2238 3872 2244 3924
rect 2052 3859 2059 3872
rect 2093 3859 2131 3872
rect 2165 3859 2203 3872
rect 2237 3859 2244 3872
rect 2052 3807 2058 3859
rect 2110 3807 2122 3859
rect 2174 3807 2186 3859
rect 2238 3807 2244 3859
rect 2052 3806 2244 3807
rect 2052 3794 2059 3806
rect 2093 3794 2131 3806
rect 2165 3794 2203 3806
rect 2237 3794 2244 3806
rect 2052 3742 2058 3794
rect 2110 3742 2122 3794
rect 2174 3742 2186 3794
rect 2238 3742 2244 3794
rect 2052 3733 2244 3742
rect 2052 3729 2059 3733
rect 2093 3729 2131 3733
rect 2165 3729 2203 3733
rect 2237 3729 2244 3733
rect 2052 3677 2058 3729
rect 2110 3677 2122 3729
rect 2174 3677 2186 3729
rect 2238 3677 2244 3729
rect 2052 3664 2244 3677
rect 2052 2972 2058 3664
rect 2238 2972 2244 3664
rect 2052 2969 2059 2972
rect 2093 2969 2131 2972
rect 2165 2969 2203 2972
rect 2237 2969 2244 2972
rect 2052 2930 2244 2969
rect 2052 2896 2059 2930
rect 2093 2896 2131 2930
rect 2165 2896 2203 2930
rect 2237 2896 2244 2930
rect 2052 2857 2244 2896
rect 2052 2823 2059 2857
rect 2093 2823 2131 2857
rect 2165 2823 2203 2857
rect 2237 2823 2244 2857
rect 2052 2784 2244 2823
rect 2052 2750 2059 2784
rect 2093 2750 2131 2784
rect 2165 2750 2203 2784
rect 2237 2750 2244 2784
rect 2052 2711 2244 2750
rect 2052 2677 2059 2711
rect 2093 2677 2131 2711
rect 2165 2677 2203 2711
rect 2237 2677 2244 2711
rect 2052 2638 2244 2677
rect 2052 2604 2059 2638
rect 2093 2604 2131 2638
rect 2165 2604 2203 2638
rect 2237 2604 2244 2638
rect 2052 2565 2244 2604
rect 2052 2531 2059 2565
rect 2093 2531 2131 2565
rect 2165 2531 2203 2565
rect 2237 2531 2244 2565
rect 2052 2492 2244 2531
rect 2052 2458 2059 2492
rect 2093 2458 2131 2492
rect 2165 2458 2203 2492
rect 2237 2458 2244 2492
rect 2052 2419 2244 2458
rect 2052 2385 2059 2419
rect 2093 2385 2131 2419
rect 2165 2385 2203 2419
rect 2237 2385 2244 2419
rect 2052 2346 2244 2385
rect 2052 2312 2059 2346
rect 2093 2312 2131 2346
rect 2165 2312 2203 2346
rect 2237 2312 2244 2346
rect 2052 2273 2244 2312
rect 2052 2239 2059 2273
rect 2093 2239 2131 2273
rect 2165 2239 2203 2273
rect 2237 2239 2244 2273
rect 2052 2200 2244 2239
rect 2052 2166 2059 2200
rect 2093 2166 2131 2200
rect 2165 2166 2203 2200
rect 2237 2166 2244 2200
rect 2052 2126 2244 2166
rect 2052 2092 2059 2126
rect 2093 2092 2131 2126
rect 2165 2092 2203 2126
rect 2237 2092 2244 2126
rect 2052 2052 2244 2092
rect 2052 2018 2059 2052
rect 2093 2018 2131 2052
rect 2165 2018 2203 2052
rect 2237 2018 2244 2052
rect 2052 1978 2244 2018
rect 2052 1944 2059 1978
rect 2093 1944 2131 1978
rect 2165 1944 2203 1978
rect 2237 1944 2244 1978
rect 2052 1904 2244 1944
rect 2052 1870 2059 1904
rect 2093 1870 2131 1904
rect 2165 1870 2203 1904
rect 2237 1870 2244 1904
rect 2052 1830 2244 1870
rect 2052 1796 2059 1830
rect 2093 1796 2131 1830
rect 2165 1796 2203 1830
rect 2237 1796 2244 1830
rect 2052 1756 2244 1796
rect 2052 1722 2059 1756
rect 2093 1722 2131 1756
rect 2165 1722 2203 1756
rect 2237 1722 2244 1756
rect 2052 1682 2244 1722
rect 2052 1648 2059 1682
rect 2093 1648 2131 1682
rect 2165 1648 2203 1682
rect 2237 1648 2244 1682
rect 2052 1608 2244 1648
rect 2052 1574 2059 1608
rect 2093 1574 2131 1608
rect 2165 1574 2203 1608
rect 2237 1574 2244 1608
rect 2052 1562 2244 1574
rect 2548 4118 2740 4130
rect 2548 4092 2627 4118
rect 2661 4092 2740 4118
rect 2548 3194 2555 4092
rect 2733 3194 2740 4092
rect 2548 3182 2740 3194
rect 2548 3148 2627 3182
rect 2661 3148 2740 3182
rect 2548 3108 2740 3148
rect 2548 3074 2555 3108
rect 2589 3074 2627 3108
rect 2661 3074 2699 3108
rect 2733 3074 2740 3108
rect 2548 3028 2740 3074
rect 2548 2994 2555 3028
rect 2589 2994 2627 3028
rect 2661 2994 2699 3028
rect 2733 2994 2740 3028
rect 2548 2948 2740 2994
rect 2548 2914 2555 2948
rect 2589 2914 2627 2948
rect 2661 2914 2699 2948
rect 2733 2914 2740 2948
rect 2548 2868 2740 2914
rect 2548 2834 2555 2868
rect 2589 2834 2627 2868
rect 2661 2834 2699 2868
rect 2733 2834 2740 2868
rect 2548 2788 2740 2834
rect 2548 2754 2555 2788
rect 2589 2754 2627 2788
rect 2661 2754 2699 2788
rect 2733 2754 2740 2788
rect 2548 2708 2740 2754
rect 2548 2674 2555 2708
rect 2589 2674 2627 2708
rect 2661 2674 2699 2708
rect 2733 2674 2740 2708
rect 2548 2657 2740 2674
rect 2548 2605 2554 2657
rect 2606 2605 2618 2657
rect 2670 2605 2682 2657
rect 2734 2605 2740 2657
rect 2548 2594 2555 2605
rect 2589 2594 2627 2605
rect 2661 2594 2699 2605
rect 2733 2594 2740 2605
rect 2548 2592 2740 2594
rect 2548 2540 2554 2592
rect 2606 2540 2618 2592
rect 2670 2540 2682 2592
rect 2734 2540 2740 2592
rect 2548 2527 2627 2540
rect 2661 2527 2740 2540
rect 2548 2475 2554 2527
rect 2606 2518 2618 2527
rect 2670 2518 2682 2527
rect 2734 2475 2740 2527
rect 2548 2462 2555 2475
rect 2733 2462 2740 2475
rect 2548 2410 2554 2462
rect 2734 2410 2740 2462
rect 2548 2397 2555 2410
rect 2733 2397 2740 2410
rect 2548 2345 2554 2397
rect 2734 2345 2740 2397
rect 2548 2332 2555 2345
rect 2733 2332 2740 2345
rect 2548 2280 2554 2332
rect 2734 2280 2740 2332
rect 2548 2267 2555 2280
rect 2733 2267 2740 2280
rect 2548 2215 2554 2267
rect 2734 2215 2740 2267
rect 2548 2202 2555 2215
rect 2733 2202 2740 2215
rect 2548 2150 2554 2202
rect 2734 2150 2740 2202
rect 2548 2137 2555 2150
rect 2733 2137 2740 2150
rect 2548 2085 2554 2137
rect 2734 2085 2740 2137
rect 2548 2072 2555 2085
rect 2733 2072 2740 2085
rect 2548 2020 2554 2072
rect 2734 2020 2740 2072
rect 2548 2007 2555 2020
rect 2733 2007 2740 2020
rect 2548 1955 2554 2007
rect 2734 1955 2740 2007
rect 2548 1942 2555 1955
rect 2733 1942 2740 1955
rect 2548 1890 2554 1942
rect 2734 1890 2740 1942
rect 2548 1877 2555 1890
rect 2733 1877 2740 1890
rect 2548 1825 2554 1877
rect 2734 1825 2740 1877
rect 2548 1812 2555 1825
rect 2733 1812 2740 1825
rect 2548 1568 2554 1812
rect 2734 1568 2740 1812
rect 2548 1562 2740 1568
rect 3044 4119 3236 4125
rect 3044 4067 3050 4119
rect 3102 4067 3114 4119
rect 3166 4067 3178 4119
rect 3230 4067 3236 4119
rect 3044 4064 3051 4067
rect 3085 4064 3123 4067
rect 3157 4064 3195 4067
rect 3229 4064 3236 4067
rect 3044 4054 3236 4064
rect 3044 4002 3050 4054
rect 3102 4002 3114 4054
rect 3166 4002 3178 4054
rect 3230 4002 3236 4054
rect 3044 3991 3051 4002
rect 3085 3991 3123 4002
rect 3157 3991 3195 4002
rect 3229 3991 3236 4002
rect 3044 3989 3236 3991
rect 3044 3937 3050 3989
rect 3102 3937 3114 3989
rect 3166 3937 3178 3989
rect 3230 3937 3236 3989
rect 3044 3924 3051 3937
rect 3085 3924 3123 3937
rect 3157 3924 3195 3937
rect 3229 3924 3236 3937
rect 3044 3872 3050 3924
rect 3102 3872 3114 3924
rect 3166 3872 3178 3924
rect 3230 3872 3236 3924
rect 3044 3859 3051 3872
rect 3085 3859 3123 3872
rect 3157 3859 3195 3872
rect 3229 3859 3236 3872
rect 3044 3807 3050 3859
rect 3102 3807 3114 3859
rect 3166 3807 3178 3859
rect 3230 3807 3236 3859
rect 3044 3806 3236 3807
rect 3044 3794 3051 3806
rect 3085 3794 3123 3806
rect 3157 3794 3195 3806
rect 3229 3794 3236 3806
rect 3044 3742 3050 3794
rect 3102 3742 3114 3794
rect 3166 3742 3178 3794
rect 3230 3742 3236 3794
rect 3044 3733 3236 3742
rect 3044 3729 3051 3733
rect 3085 3729 3123 3733
rect 3157 3729 3195 3733
rect 3229 3729 3236 3733
rect 3044 3677 3050 3729
rect 3102 3677 3114 3729
rect 3166 3677 3178 3729
rect 3230 3677 3236 3729
rect 3044 3664 3236 3677
rect 3044 2972 3050 3664
rect 3230 2972 3236 3664
rect 3044 2969 3051 2972
rect 3085 2969 3123 2972
rect 3157 2969 3195 2972
rect 3229 2969 3236 2972
rect 3044 2930 3236 2969
rect 3044 2896 3051 2930
rect 3085 2896 3123 2930
rect 3157 2896 3195 2930
rect 3229 2896 3236 2930
rect 3044 2857 3236 2896
rect 3044 2823 3051 2857
rect 3085 2823 3123 2857
rect 3157 2823 3195 2857
rect 3229 2823 3236 2857
rect 3044 2784 3236 2823
rect 3044 2750 3051 2784
rect 3085 2750 3123 2784
rect 3157 2750 3195 2784
rect 3229 2750 3236 2784
rect 3044 2711 3236 2750
rect 3044 2677 3051 2711
rect 3085 2677 3123 2711
rect 3157 2677 3195 2711
rect 3229 2677 3236 2711
rect 3044 2638 3236 2677
rect 3044 2604 3051 2638
rect 3085 2604 3123 2638
rect 3157 2604 3195 2638
rect 3229 2604 3236 2638
rect 3044 2565 3236 2604
rect 3044 2531 3051 2565
rect 3085 2531 3123 2565
rect 3157 2531 3195 2565
rect 3229 2531 3236 2565
rect 3044 2492 3236 2531
rect 3044 2458 3051 2492
rect 3085 2458 3123 2492
rect 3157 2458 3195 2492
rect 3229 2458 3236 2492
rect 3044 2419 3236 2458
rect 3044 2385 3051 2419
rect 3085 2385 3123 2419
rect 3157 2385 3195 2419
rect 3229 2385 3236 2419
rect 3044 2346 3236 2385
rect 3044 2312 3051 2346
rect 3085 2312 3123 2346
rect 3157 2312 3195 2346
rect 3229 2312 3236 2346
rect 3044 2273 3236 2312
rect 3044 2239 3051 2273
rect 3085 2239 3123 2273
rect 3157 2239 3195 2273
rect 3229 2239 3236 2273
rect 3044 2200 3236 2239
rect 3044 2166 3051 2200
rect 3085 2166 3123 2200
rect 3157 2166 3195 2200
rect 3229 2166 3236 2200
rect 3044 2126 3236 2166
rect 3044 2092 3051 2126
rect 3085 2092 3123 2126
rect 3157 2092 3195 2126
rect 3229 2092 3236 2126
rect 3044 2052 3236 2092
rect 3044 2018 3051 2052
rect 3085 2018 3123 2052
rect 3157 2018 3195 2052
rect 3229 2018 3236 2052
rect 3044 1978 3236 2018
rect 3044 1944 3051 1978
rect 3085 1944 3123 1978
rect 3157 1944 3195 1978
rect 3229 1944 3236 1978
rect 3044 1904 3236 1944
rect 3044 1870 3051 1904
rect 3085 1870 3123 1904
rect 3157 1870 3195 1904
rect 3229 1870 3236 1904
rect 3044 1830 3236 1870
rect 3044 1796 3051 1830
rect 3085 1796 3123 1830
rect 3157 1796 3195 1830
rect 3229 1796 3236 1830
rect 3044 1756 3236 1796
rect 3044 1722 3051 1756
rect 3085 1722 3123 1756
rect 3157 1722 3195 1756
rect 3229 1722 3236 1756
rect 3044 1682 3236 1722
rect 3044 1648 3051 1682
rect 3085 1648 3123 1682
rect 3157 1648 3195 1682
rect 3229 1648 3236 1682
rect 3044 1608 3236 1648
rect 3044 1574 3051 1608
rect 3085 1574 3123 1608
rect 3157 1574 3195 1608
rect 3229 1574 3236 1608
rect 3044 1562 3236 1574
rect 3540 4118 3732 4130
rect 3540 4092 3619 4118
rect 3653 4092 3732 4118
rect 3540 3194 3547 4092
rect 3725 3194 3732 4092
rect 3540 3182 3732 3194
rect 3540 3148 3619 3182
rect 3653 3148 3732 3182
rect 3540 3108 3732 3148
rect 3540 3074 3547 3108
rect 3581 3074 3619 3108
rect 3653 3074 3691 3108
rect 3725 3074 3732 3108
rect 3540 3028 3732 3074
rect 3540 2994 3547 3028
rect 3581 2994 3619 3028
rect 3653 2994 3691 3028
rect 3725 2994 3732 3028
rect 3540 2948 3732 2994
rect 3540 2914 3547 2948
rect 3581 2914 3619 2948
rect 3653 2914 3691 2948
rect 3725 2914 3732 2948
rect 3540 2868 3732 2914
rect 3540 2834 3547 2868
rect 3581 2834 3619 2868
rect 3653 2834 3691 2868
rect 3725 2834 3732 2868
rect 3540 2788 3732 2834
rect 3540 2754 3547 2788
rect 3581 2754 3619 2788
rect 3653 2754 3691 2788
rect 3725 2754 3732 2788
rect 3540 2708 3732 2754
rect 3540 2674 3547 2708
rect 3581 2674 3619 2708
rect 3653 2674 3691 2708
rect 3725 2674 3732 2708
rect 3540 2657 3732 2674
rect 3540 2605 3546 2657
rect 3598 2605 3610 2657
rect 3662 2605 3674 2657
rect 3726 2605 3732 2657
rect 3540 2594 3547 2605
rect 3581 2594 3619 2605
rect 3653 2594 3691 2605
rect 3725 2594 3732 2605
rect 3540 2592 3732 2594
rect 3540 2540 3546 2592
rect 3598 2540 3610 2592
rect 3662 2540 3674 2592
rect 3726 2540 3732 2592
rect 3540 2527 3619 2540
rect 3653 2527 3732 2540
rect 3540 2475 3546 2527
rect 3598 2518 3610 2527
rect 3662 2518 3674 2527
rect 3726 2475 3732 2527
rect 3540 2462 3547 2475
rect 3725 2462 3732 2475
rect 3540 2410 3546 2462
rect 3726 2410 3732 2462
rect 3540 2397 3547 2410
rect 3725 2397 3732 2410
rect 3540 2345 3546 2397
rect 3726 2345 3732 2397
rect 3540 2332 3547 2345
rect 3725 2332 3732 2345
rect 3540 2280 3546 2332
rect 3726 2280 3732 2332
rect 3540 2267 3547 2280
rect 3725 2267 3732 2280
rect 3540 2215 3546 2267
rect 3726 2215 3732 2267
rect 3540 2202 3547 2215
rect 3725 2202 3732 2215
rect 3540 2150 3546 2202
rect 3726 2150 3732 2202
rect 3540 2137 3547 2150
rect 3725 2137 3732 2150
rect 3540 2085 3546 2137
rect 3726 2085 3732 2137
rect 3540 2072 3547 2085
rect 3725 2072 3732 2085
rect 3540 2020 3546 2072
rect 3726 2020 3732 2072
rect 3540 2007 3547 2020
rect 3725 2007 3732 2020
rect 3540 1955 3546 2007
rect 3726 1955 3732 2007
rect 3540 1942 3547 1955
rect 3725 1942 3732 1955
rect 3540 1890 3546 1942
rect 3726 1890 3732 1942
rect 3540 1877 3547 1890
rect 3725 1877 3732 1890
rect 3540 1825 3546 1877
rect 3726 1825 3732 1877
rect 3540 1812 3547 1825
rect 3725 1812 3732 1825
rect 3540 1568 3546 1812
rect 3726 1568 3732 1812
rect 3540 1562 3732 1568
rect 4036 4119 4228 4125
rect 4036 4067 4042 4119
rect 4094 4067 4106 4119
rect 4158 4067 4170 4119
rect 4222 4067 4228 4119
rect 4036 4064 4043 4067
rect 4077 4064 4115 4067
rect 4149 4064 4187 4067
rect 4221 4064 4228 4067
rect 4036 4054 4228 4064
rect 4036 4002 4042 4054
rect 4094 4002 4106 4054
rect 4158 4002 4170 4054
rect 4222 4002 4228 4054
rect 4036 3991 4043 4002
rect 4077 3991 4115 4002
rect 4149 3991 4187 4002
rect 4221 3991 4228 4002
rect 4036 3989 4228 3991
rect 4036 3937 4042 3989
rect 4094 3937 4106 3989
rect 4158 3937 4170 3989
rect 4222 3937 4228 3989
rect 4036 3924 4043 3937
rect 4077 3924 4115 3937
rect 4149 3924 4187 3937
rect 4221 3924 4228 3937
rect 4036 3872 4042 3924
rect 4094 3872 4106 3924
rect 4158 3872 4170 3924
rect 4222 3872 4228 3924
rect 4036 3859 4043 3872
rect 4077 3859 4115 3872
rect 4149 3859 4187 3872
rect 4221 3859 4228 3872
rect 4036 3807 4042 3859
rect 4094 3807 4106 3859
rect 4158 3807 4170 3859
rect 4222 3807 4228 3859
rect 4036 3806 4228 3807
rect 4036 3794 4043 3806
rect 4077 3794 4115 3806
rect 4149 3794 4187 3806
rect 4221 3794 4228 3806
rect 4036 3742 4042 3794
rect 4094 3742 4106 3794
rect 4158 3742 4170 3794
rect 4222 3742 4228 3794
rect 4036 3733 4228 3742
rect 4036 3729 4043 3733
rect 4077 3729 4115 3733
rect 4149 3729 4187 3733
rect 4221 3729 4228 3733
rect 4036 3677 4042 3729
rect 4094 3677 4106 3729
rect 4158 3677 4170 3729
rect 4222 3677 4228 3729
rect 4036 3664 4228 3677
rect 4036 2972 4042 3664
rect 4222 2972 4228 3664
rect 4036 2969 4043 2972
rect 4077 2969 4115 2972
rect 4149 2969 4187 2972
rect 4221 2969 4228 2972
rect 4036 2930 4228 2969
rect 4036 2896 4043 2930
rect 4077 2896 4115 2930
rect 4149 2896 4187 2930
rect 4221 2896 4228 2930
rect 4036 2857 4228 2896
rect 4036 2823 4043 2857
rect 4077 2823 4115 2857
rect 4149 2823 4187 2857
rect 4221 2823 4228 2857
rect 4036 2784 4228 2823
rect 4036 2750 4043 2784
rect 4077 2750 4115 2784
rect 4149 2750 4187 2784
rect 4221 2750 4228 2784
rect 4036 2711 4228 2750
rect 4036 2677 4043 2711
rect 4077 2677 4115 2711
rect 4149 2677 4187 2711
rect 4221 2677 4228 2711
rect 4036 2638 4228 2677
rect 4036 2604 4043 2638
rect 4077 2604 4115 2638
rect 4149 2604 4187 2638
rect 4221 2604 4228 2638
rect 4036 2565 4228 2604
rect 4036 2531 4043 2565
rect 4077 2531 4115 2565
rect 4149 2531 4187 2565
rect 4221 2531 4228 2565
rect 4036 2492 4228 2531
rect 4036 2458 4043 2492
rect 4077 2458 4115 2492
rect 4149 2458 4187 2492
rect 4221 2458 4228 2492
rect 4036 2419 4228 2458
rect 4036 2385 4043 2419
rect 4077 2385 4115 2419
rect 4149 2385 4187 2419
rect 4221 2385 4228 2419
rect 4036 2346 4228 2385
rect 4036 2312 4043 2346
rect 4077 2312 4115 2346
rect 4149 2312 4187 2346
rect 4221 2312 4228 2346
rect 4036 2273 4228 2312
rect 4036 2239 4043 2273
rect 4077 2239 4115 2273
rect 4149 2239 4187 2273
rect 4221 2239 4228 2273
rect 4036 2200 4228 2239
rect 4036 2166 4043 2200
rect 4077 2166 4115 2200
rect 4149 2166 4187 2200
rect 4221 2166 4228 2200
rect 4036 2126 4228 2166
rect 4036 2092 4043 2126
rect 4077 2092 4115 2126
rect 4149 2092 4187 2126
rect 4221 2092 4228 2126
rect 4036 2052 4228 2092
rect 4036 2018 4043 2052
rect 4077 2018 4115 2052
rect 4149 2018 4187 2052
rect 4221 2018 4228 2052
rect 4036 1978 4228 2018
rect 4036 1944 4043 1978
rect 4077 1944 4115 1978
rect 4149 1944 4187 1978
rect 4221 1944 4228 1978
rect 4036 1904 4228 1944
rect 4036 1870 4043 1904
rect 4077 1870 4115 1904
rect 4149 1870 4187 1904
rect 4221 1870 4228 1904
rect 4036 1830 4228 1870
rect 4036 1796 4043 1830
rect 4077 1796 4115 1830
rect 4149 1796 4187 1830
rect 4221 1796 4228 1830
rect 4036 1756 4228 1796
rect 4036 1722 4043 1756
rect 4077 1722 4115 1756
rect 4149 1722 4187 1756
rect 4221 1722 4228 1756
rect 4036 1682 4228 1722
rect 4036 1648 4043 1682
rect 4077 1648 4115 1682
rect 4149 1648 4187 1682
rect 4221 1648 4228 1682
rect 4036 1608 4228 1648
rect 4036 1574 4043 1608
rect 4077 1574 4115 1608
rect 4149 1574 4187 1608
rect 4221 1574 4228 1608
rect 4036 1562 4228 1574
rect 4532 4118 4724 4130
rect 4532 4092 4611 4118
rect 4645 4092 4724 4118
rect 4532 3194 4539 4092
rect 4717 3194 4724 4092
rect 4532 3182 4724 3194
rect 4532 3148 4611 3182
rect 4645 3148 4724 3182
rect 4532 3108 4724 3148
rect 4532 3074 4539 3108
rect 4573 3074 4611 3108
rect 4645 3074 4683 3108
rect 4717 3074 4724 3108
rect 4532 3028 4724 3074
rect 4532 2994 4539 3028
rect 4573 2994 4611 3028
rect 4645 2994 4683 3028
rect 4717 2994 4724 3028
rect 4532 2948 4724 2994
rect 4532 2914 4539 2948
rect 4573 2914 4611 2948
rect 4645 2914 4683 2948
rect 4717 2914 4724 2948
rect 4532 2868 4724 2914
rect 4532 2834 4539 2868
rect 4573 2834 4611 2868
rect 4645 2834 4683 2868
rect 4717 2834 4724 2868
rect 4532 2788 4724 2834
rect 4532 2754 4539 2788
rect 4573 2754 4611 2788
rect 4645 2754 4683 2788
rect 4717 2754 4724 2788
rect 4532 2708 4724 2754
rect 4532 2674 4539 2708
rect 4573 2674 4611 2708
rect 4645 2674 4683 2708
rect 4717 2674 4724 2708
rect 4532 2657 4724 2674
rect 4532 2605 4538 2657
rect 4590 2605 4602 2657
rect 4654 2605 4666 2657
rect 4718 2605 4724 2657
rect 4532 2594 4539 2605
rect 4573 2594 4611 2605
rect 4645 2594 4683 2605
rect 4717 2594 4724 2605
rect 4532 2592 4724 2594
rect 4532 2540 4538 2592
rect 4590 2540 4602 2592
rect 4654 2540 4666 2592
rect 4718 2540 4724 2592
rect 4532 2527 4611 2540
rect 4645 2527 4724 2540
rect 4532 2475 4538 2527
rect 4590 2518 4602 2527
rect 4654 2518 4666 2527
rect 4718 2475 4724 2527
rect 4532 2462 4539 2475
rect 4717 2462 4724 2475
rect 4532 2410 4538 2462
rect 4718 2410 4724 2462
rect 4532 2397 4539 2410
rect 4717 2397 4724 2410
rect 4532 2345 4538 2397
rect 4718 2345 4724 2397
rect 4532 2332 4539 2345
rect 4717 2332 4724 2345
rect 4532 2280 4538 2332
rect 4718 2280 4724 2332
rect 4532 2267 4539 2280
rect 4717 2267 4724 2280
rect 4532 2215 4538 2267
rect 4718 2215 4724 2267
rect 4532 2202 4539 2215
rect 4717 2202 4724 2215
rect 4532 2150 4538 2202
rect 4718 2150 4724 2202
rect 4532 2137 4539 2150
rect 4717 2137 4724 2150
rect 4532 2085 4538 2137
rect 4718 2085 4724 2137
rect 4532 2072 4539 2085
rect 4717 2072 4724 2085
rect 4532 2020 4538 2072
rect 4718 2020 4724 2072
rect 4532 2007 4539 2020
rect 4717 2007 4724 2020
rect 4532 1955 4538 2007
rect 4718 1955 4724 2007
rect 4532 1942 4539 1955
rect 4717 1942 4724 1955
rect 4532 1890 4538 1942
rect 4718 1890 4724 1942
rect 4532 1877 4539 1890
rect 4717 1877 4724 1890
rect 4532 1825 4538 1877
rect 4718 1825 4724 1877
rect 4532 1812 4539 1825
rect 4717 1812 4724 1825
rect 4532 1568 4538 1812
rect 4718 1568 4724 1812
rect 4532 1562 4724 1568
rect 5028 4119 5220 4125
rect 5028 4067 5034 4119
rect 5086 4067 5098 4119
rect 5150 4067 5162 4119
rect 5214 4067 5220 4119
rect 5028 4064 5035 4067
rect 5069 4064 5107 4067
rect 5141 4064 5179 4067
rect 5213 4064 5220 4067
rect 5028 4054 5220 4064
rect 5028 4002 5034 4054
rect 5086 4002 5098 4054
rect 5150 4002 5162 4054
rect 5214 4002 5220 4054
rect 5028 3991 5035 4002
rect 5069 3991 5107 4002
rect 5141 3991 5179 4002
rect 5213 3991 5220 4002
rect 5028 3989 5220 3991
rect 5028 3937 5034 3989
rect 5086 3937 5098 3989
rect 5150 3937 5162 3989
rect 5214 3937 5220 3989
rect 5028 3924 5035 3937
rect 5069 3924 5107 3937
rect 5141 3924 5179 3937
rect 5213 3924 5220 3937
rect 5028 3872 5034 3924
rect 5086 3872 5098 3924
rect 5150 3872 5162 3924
rect 5214 3872 5220 3924
rect 5028 3859 5035 3872
rect 5069 3859 5107 3872
rect 5141 3859 5179 3872
rect 5213 3859 5220 3872
rect 5028 3807 5034 3859
rect 5086 3807 5098 3859
rect 5150 3807 5162 3859
rect 5214 3807 5220 3859
rect 5028 3806 5220 3807
rect 5028 3794 5035 3806
rect 5069 3794 5107 3806
rect 5141 3794 5179 3806
rect 5213 3794 5220 3806
rect 5028 3742 5034 3794
rect 5086 3742 5098 3794
rect 5150 3742 5162 3794
rect 5214 3742 5220 3794
rect 5028 3733 5220 3742
rect 5028 3729 5035 3733
rect 5069 3729 5107 3733
rect 5141 3729 5179 3733
rect 5213 3729 5220 3733
rect 5028 3677 5034 3729
rect 5086 3677 5098 3729
rect 5150 3677 5162 3729
rect 5214 3677 5220 3729
rect 5028 3664 5220 3677
rect 5028 2972 5034 3664
rect 5214 2972 5220 3664
rect 5028 2969 5035 2972
rect 5069 2969 5107 2972
rect 5141 2969 5179 2972
rect 5213 2969 5220 2972
rect 5028 2930 5220 2969
rect 5028 2896 5035 2930
rect 5069 2896 5107 2930
rect 5141 2896 5179 2930
rect 5213 2896 5220 2930
rect 5028 2857 5220 2896
rect 5028 2823 5035 2857
rect 5069 2823 5107 2857
rect 5141 2823 5179 2857
rect 5213 2823 5220 2857
rect 5028 2784 5220 2823
rect 5028 2750 5035 2784
rect 5069 2750 5107 2784
rect 5141 2750 5179 2784
rect 5213 2750 5220 2784
rect 5028 2711 5220 2750
rect 5028 2677 5035 2711
rect 5069 2677 5107 2711
rect 5141 2677 5179 2711
rect 5213 2677 5220 2711
rect 5028 2638 5220 2677
rect 5028 2604 5035 2638
rect 5069 2604 5107 2638
rect 5141 2604 5179 2638
rect 5213 2604 5220 2638
rect 5028 2565 5220 2604
rect 5028 2531 5035 2565
rect 5069 2531 5107 2565
rect 5141 2531 5179 2565
rect 5213 2531 5220 2565
rect 5028 2492 5220 2531
rect 5028 2458 5035 2492
rect 5069 2458 5107 2492
rect 5141 2458 5179 2492
rect 5213 2458 5220 2492
rect 5028 2419 5220 2458
rect 5028 2385 5035 2419
rect 5069 2385 5107 2419
rect 5141 2385 5179 2419
rect 5213 2385 5220 2419
rect 5028 2346 5220 2385
rect 5028 2312 5035 2346
rect 5069 2312 5107 2346
rect 5141 2312 5179 2346
rect 5213 2312 5220 2346
rect 5028 2273 5220 2312
rect 5028 2239 5035 2273
rect 5069 2239 5107 2273
rect 5141 2239 5179 2273
rect 5213 2239 5220 2273
rect 5028 2200 5220 2239
rect 5028 2166 5035 2200
rect 5069 2166 5107 2200
rect 5141 2166 5179 2200
rect 5213 2166 5220 2200
rect 5028 2126 5220 2166
rect 5028 2092 5035 2126
rect 5069 2092 5107 2126
rect 5141 2092 5179 2126
rect 5213 2092 5220 2126
rect 5028 2052 5220 2092
rect 5028 2018 5035 2052
rect 5069 2018 5107 2052
rect 5141 2018 5179 2052
rect 5213 2018 5220 2052
rect 5028 1978 5220 2018
rect 5028 1944 5035 1978
rect 5069 1944 5107 1978
rect 5141 1944 5179 1978
rect 5213 1944 5220 1978
rect 5028 1904 5220 1944
rect 5028 1870 5035 1904
rect 5069 1870 5107 1904
rect 5141 1870 5179 1904
rect 5213 1870 5220 1904
rect 5028 1830 5220 1870
rect 5028 1796 5035 1830
rect 5069 1796 5107 1830
rect 5141 1796 5179 1830
rect 5213 1796 5220 1830
rect 5028 1756 5220 1796
rect 5028 1722 5035 1756
rect 5069 1722 5107 1756
rect 5141 1722 5179 1756
rect 5213 1722 5220 1756
rect 5028 1682 5220 1722
rect 5028 1648 5035 1682
rect 5069 1648 5107 1682
rect 5141 1648 5179 1682
rect 5213 1648 5220 1682
rect 5028 1608 5220 1648
rect 5028 1574 5035 1608
rect 5069 1574 5107 1608
rect 5141 1574 5179 1608
rect 5213 1574 5220 1608
rect 5028 1562 5220 1574
rect 5524 4118 5716 4130
rect 5524 4092 5603 4118
rect 5637 4092 5716 4118
rect 5524 3194 5531 4092
rect 5709 3194 5716 4092
rect 5524 3182 5716 3194
rect 5524 3148 5603 3182
rect 5637 3148 5716 3182
rect 5524 3108 5716 3148
rect 5524 3074 5531 3108
rect 5565 3074 5603 3108
rect 5637 3074 5675 3108
rect 5709 3074 5716 3108
rect 5524 3028 5716 3074
rect 5524 2994 5531 3028
rect 5565 2994 5603 3028
rect 5637 2994 5675 3028
rect 5709 2994 5716 3028
rect 5524 2948 5716 2994
rect 5524 2914 5531 2948
rect 5565 2914 5603 2948
rect 5637 2914 5675 2948
rect 5709 2914 5716 2948
rect 5524 2868 5716 2914
rect 5524 2834 5531 2868
rect 5565 2834 5603 2868
rect 5637 2834 5675 2868
rect 5709 2834 5716 2868
rect 5524 2788 5716 2834
rect 5524 2754 5531 2788
rect 5565 2754 5603 2788
rect 5637 2754 5675 2788
rect 5709 2754 5716 2788
rect 5524 2708 5716 2754
rect 5524 2674 5531 2708
rect 5565 2674 5603 2708
rect 5637 2674 5675 2708
rect 5709 2674 5716 2708
rect 5524 2657 5716 2674
rect 5524 2605 5530 2657
rect 5582 2605 5594 2657
rect 5646 2605 5658 2657
rect 5710 2605 5716 2657
rect 5524 2594 5531 2605
rect 5565 2594 5603 2605
rect 5637 2594 5675 2605
rect 5709 2594 5716 2605
rect 5524 2592 5716 2594
rect 5524 2540 5530 2592
rect 5582 2540 5594 2592
rect 5646 2540 5658 2592
rect 5710 2540 5716 2592
rect 5524 2527 5603 2540
rect 5637 2527 5716 2540
rect 5524 2475 5530 2527
rect 5582 2518 5594 2527
rect 5646 2518 5658 2527
rect 5710 2475 5716 2527
rect 5524 2462 5531 2475
rect 5709 2462 5716 2475
rect 5524 2410 5530 2462
rect 5710 2410 5716 2462
rect 5524 2397 5531 2410
rect 5709 2397 5716 2410
rect 5524 2345 5530 2397
rect 5710 2345 5716 2397
rect 5524 2332 5531 2345
rect 5709 2332 5716 2345
rect 5524 2280 5530 2332
rect 5710 2280 5716 2332
rect 5524 2267 5531 2280
rect 5709 2267 5716 2280
rect 5524 2215 5530 2267
rect 5710 2215 5716 2267
rect 5524 2202 5531 2215
rect 5709 2202 5716 2215
rect 5524 2150 5530 2202
rect 5710 2150 5716 2202
rect 5524 2137 5531 2150
rect 5709 2137 5716 2150
rect 5524 2085 5530 2137
rect 5710 2085 5716 2137
rect 5524 2072 5531 2085
rect 5709 2072 5716 2085
rect 5524 2020 5530 2072
rect 5710 2020 5716 2072
rect 5524 2007 5531 2020
rect 5709 2007 5716 2020
rect 5524 1955 5530 2007
rect 5710 1955 5716 2007
rect 5524 1942 5531 1955
rect 5709 1942 5716 1955
rect 5524 1890 5530 1942
rect 5710 1890 5716 1942
rect 5524 1877 5531 1890
rect 5709 1877 5716 1890
rect 5524 1825 5530 1877
rect 5710 1825 5716 1877
rect 5524 1812 5531 1825
rect 5709 1812 5716 1825
rect 5524 1568 5530 1812
rect 5710 1568 5716 1812
rect 5524 1562 5716 1568
rect 6020 4119 6212 4125
rect 6020 4067 6026 4119
rect 6078 4067 6090 4119
rect 6142 4067 6154 4119
rect 6206 4067 6212 4119
rect 6020 4064 6027 4067
rect 6061 4064 6099 4067
rect 6133 4064 6171 4067
rect 6205 4064 6212 4067
rect 6020 4054 6212 4064
rect 6020 4002 6026 4054
rect 6078 4002 6090 4054
rect 6142 4002 6154 4054
rect 6206 4002 6212 4054
rect 6020 3991 6027 4002
rect 6061 3991 6099 4002
rect 6133 3991 6171 4002
rect 6205 3991 6212 4002
rect 6020 3989 6212 3991
rect 6020 3937 6026 3989
rect 6078 3937 6090 3989
rect 6142 3937 6154 3989
rect 6206 3937 6212 3989
rect 6020 3924 6027 3937
rect 6061 3924 6099 3937
rect 6133 3924 6171 3937
rect 6205 3924 6212 3937
rect 6020 3872 6026 3924
rect 6078 3872 6090 3924
rect 6142 3872 6154 3924
rect 6206 3872 6212 3924
rect 6020 3859 6027 3872
rect 6061 3859 6099 3872
rect 6133 3859 6171 3872
rect 6205 3859 6212 3872
rect 6020 3807 6026 3859
rect 6078 3807 6090 3859
rect 6142 3807 6154 3859
rect 6206 3807 6212 3859
rect 6020 3806 6212 3807
rect 6020 3794 6027 3806
rect 6061 3794 6099 3806
rect 6133 3794 6171 3806
rect 6205 3794 6212 3806
rect 6020 3742 6026 3794
rect 6078 3742 6090 3794
rect 6142 3742 6154 3794
rect 6206 3742 6212 3794
rect 6020 3733 6212 3742
rect 6020 3729 6027 3733
rect 6061 3729 6099 3733
rect 6133 3729 6171 3733
rect 6205 3729 6212 3733
rect 6020 3677 6026 3729
rect 6078 3677 6090 3729
rect 6142 3677 6154 3729
rect 6206 3677 6212 3729
rect 6020 3664 6212 3677
rect 6020 2972 6026 3664
rect 6206 2972 6212 3664
rect 6020 2969 6027 2972
rect 6061 2969 6099 2972
rect 6133 2969 6171 2972
rect 6205 2969 6212 2972
rect 6020 2930 6212 2969
rect 6020 2896 6027 2930
rect 6061 2896 6099 2930
rect 6133 2896 6171 2930
rect 6205 2896 6212 2930
rect 6020 2857 6212 2896
rect 6020 2823 6027 2857
rect 6061 2823 6099 2857
rect 6133 2823 6171 2857
rect 6205 2823 6212 2857
rect 6020 2784 6212 2823
rect 6020 2750 6027 2784
rect 6061 2750 6099 2784
rect 6133 2750 6171 2784
rect 6205 2750 6212 2784
rect 6020 2711 6212 2750
rect 6020 2677 6027 2711
rect 6061 2677 6099 2711
rect 6133 2677 6171 2711
rect 6205 2677 6212 2711
rect 6020 2638 6212 2677
rect 6020 2604 6027 2638
rect 6061 2604 6099 2638
rect 6133 2604 6171 2638
rect 6205 2604 6212 2638
rect 6020 2565 6212 2604
rect 6020 2531 6027 2565
rect 6061 2531 6099 2565
rect 6133 2531 6171 2565
rect 6205 2531 6212 2565
rect 6020 2492 6212 2531
rect 6020 2458 6027 2492
rect 6061 2458 6099 2492
rect 6133 2458 6171 2492
rect 6205 2458 6212 2492
rect 6020 2419 6212 2458
rect 6020 2385 6027 2419
rect 6061 2385 6099 2419
rect 6133 2385 6171 2419
rect 6205 2385 6212 2419
rect 6020 2346 6212 2385
rect 6020 2312 6027 2346
rect 6061 2312 6099 2346
rect 6133 2312 6171 2346
rect 6205 2312 6212 2346
rect 6020 2273 6212 2312
rect 6020 2239 6027 2273
rect 6061 2239 6099 2273
rect 6133 2239 6171 2273
rect 6205 2239 6212 2273
rect 6020 2200 6212 2239
rect 6020 2166 6027 2200
rect 6061 2166 6099 2200
rect 6133 2166 6171 2200
rect 6205 2166 6212 2200
rect 6020 2126 6212 2166
rect 6020 2092 6027 2126
rect 6061 2092 6099 2126
rect 6133 2092 6171 2126
rect 6205 2092 6212 2126
rect 6020 2052 6212 2092
rect 6020 2018 6027 2052
rect 6061 2018 6099 2052
rect 6133 2018 6171 2052
rect 6205 2018 6212 2052
rect 6020 1978 6212 2018
rect 6020 1944 6027 1978
rect 6061 1944 6099 1978
rect 6133 1944 6171 1978
rect 6205 1944 6212 1978
rect 6020 1904 6212 1944
rect 6020 1870 6027 1904
rect 6061 1870 6099 1904
rect 6133 1870 6171 1904
rect 6205 1870 6212 1904
rect 6020 1830 6212 1870
rect 6020 1796 6027 1830
rect 6061 1796 6099 1830
rect 6133 1796 6171 1830
rect 6205 1796 6212 1830
rect 6020 1756 6212 1796
rect 6020 1722 6027 1756
rect 6061 1722 6099 1756
rect 6133 1722 6171 1756
rect 6205 1722 6212 1756
rect 6020 1682 6212 1722
rect 6020 1648 6027 1682
rect 6061 1648 6099 1682
rect 6133 1648 6171 1682
rect 6205 1648 6212 1682
rect 6020 1608 6212 1648
rect 6020 1574 6027 1608
rect 6061 1574 6099 1608
rect 6133 1574 6171 1608
rect 6205 1574 6212 1608
rect 6020 1562 6212 1574
rect 6516 4118 6708 4130
rect 6516 4092 6595 4118
rect 6629 4092 6708 4118
rect 6516 3194 6523 4092
rect 6701 3194 6708 4092
rect 6516 3182 6708 3194
rect 6516 3148 6595 3182
rect 6629 3148 6708 3182
rect 6516 3108 6708 3148
rect 6516 3074 6523 3108
rect 6557 3074 6595 3108
rect 6629 3074 6667 3108
rect 6701 3074 6708 3108
rect 6516 3028 6708 3074
rect 6516 2994 6523 3028
rect 6557 2994 6595 3028
rect 6629 2994 6667 3028
rect 6701 2994 6708 3028
rect 6516 2948 6708 2994
rect 6516 2914 6523 2948
rect 6557 2914 6595 2948
rect 6629 2914 6667 2948
rect 6701 2914 6708 2948
rect 6516 2868 6708 2914
rect 6516 2834 6523 2868
rect 6557 2834 6595 2868
rect 6629 2834 6667 2868
rect 6701 2834 6708 2868
rect 6516 2788 6708 2834
rect 6516 2754 6523 2788
rect 6557 2754 6595 2788
rect 6629 2754 6667 2788
rect 6701 2754 6708 2788
rect 6516 2708 6708 2754
rect 6516 2674 6523 2708
rect 6557 2674 6595 2708
rect 6629 2674 6667 2708
rect 6701 2674 6708 2708
rect 6516 2657 6708 2674
rect 6516 2605 6522 2657
rect 6574 2605 6586 2657
rect 6638 2605 6650 2657
rect 6702 2605 6708 2657
rect 6516 2594 6523 2605
rect 6557 2594 6595 2605
rect 6629 2594 6667 2605
rect 6701 2594 6708 2605
rect 6516 2592 6708 2594
rect 6516 2540 6522 2592
rect 6574 2540 6586 2592
rect 6638 2540 6650 2592
rect 6702 2540 6708 2592
rect 6516 2527 6595 2540
rect 6629 2527 6708 2540
rect 6516 2475 6522 2527
rect 6574 2518 6586 2527
rect 6638 2518 6650 2527
rect 6702 2475 6708 2527
rect 6516 2462 6523 2475
rect 6701 2462 6708 2475
rect 6516 2410 6522 2462
rect 6702 2410 6708 2462
rect 6516 2397 6523 2410
rect 6701 2397 6708 2410
rect 6516 2345 6522 2397
rect 6702 2345 6708 2397
rect 6516 2332 6523 2345
rect 6701 2332 6708 2345
rect 6516 2280 6522 2332
rect 6702 2280 6708 2332
rect 6516 2267 6523 2280
rect 6701 2267 6708 2280
rect 6516 2215 6522 2267
rect 6702 2215 6708 2267
rect 6516 2202 6523 2215
rect 6701 2202 6708 2215
rect 6516 2150 6522 2202
rect 6702 2150 6708 2202
rect 6516 2137 6523 2150
rect 6701 2137 6708 2150
rect 6516 2085 6522 2137
rect 6702 2085 6708 2137
rect 6516 2072 6523 2085
rect 6701 2072 6708 2085
rect 6516 2020 6522 2072
rect 6702 2020 6708 2072
rect 6516 2007 6523 2020
rect 6701 2007 6708 2020
rect 6516 1955 6522 2007
rect 6702 1955 6708 2007
rect 6516 1942 6523 1955
rect 6701 1942 6708 1955
rect 6516 1890 6522 1942
rect 6702 1890 6708 1942
rect 6516 1877 6523 1890
rect 6701 1877 6708 1890
rect 6516 1825 6522 1877
rect 6702 1825 6708 1877
rect 6516 1812 6523 1825
rect 6701 1812 6708 1825
rect 6516 1568 6522 1812
rect 6702 1568 6708 1812
rect 6516 1562 6708 1568
rect 7012 4119 7204 4125
rect 7012 4067 7018 4119
rect 7070 4067 7082 4119
rect 7134 4067 7146 4119
rect 7198 4067 7204 4119
rect 7012 4064 7019 4067
rect 7053 4064 7091 4067
rect 7125 4064 7163 4067
rect 7197 4064 7204 4067
rect 7012 4054 7204 4064
rect 7012 4002 7018 4054
rect 7070 4002 7082 4054
rect 7134 4002 7146 4054
rect 7198 4002 7204 4054
rect 7012 3991 7019 4002
rect 7053 3991 7091 4002
rect 7125 3991 7163 4002
rect 7197 3991 7204 4002
rect 7012 3989 7204 3991
rect 7012 3937 7018 3989
rect 7070 3937 7082 3989
rect 7134 3937 7146 3989
rect 7198 3937 7204 3989
rect 7012 3924 7019 3937
rect 7053 3924 7091 3937
rect 7125 3924 7163 3937
rect 7197 3924 7204 3937
rect 7012 3872 7018 3924
rect 7070 3872 7082 3924
rect 7134 3872 7146 3924
rect 7198 3872 7204 3924
rect 7012 3859 7019 3872
rect 7053 3859 7091 3872
rect 7125 3859 7163 3872
rect 7197 3859 7204 3872
rect 7012 3807 7018 3859
rect 7070 3807 7082 3859
rect 7134 3807 7146 3859
rect 7198 3807 7204 3859
rect 7012 3806 7204 3807
rect 7012 3794 7019 3806
rect 7053 3794 7091 3806
rect 7125 3794 7163 3806
rect 7197 3794 7204 3806
rect 7012 3742 7018 3794
rect 7070 3742 7082 3794
rect 7134 3742 7146 3794
rect 7198 3742 7204 3794
rect 7012 3733 7204 3742
rect 7012 3729 7019 3733
rect 7053 3729 7091 3733
rect 7125 3729 7163 3733
rect 7197 3729 7204 3733
rect 7012 3677 7018 3729
rect 7070 3677 7082 3729
rect 7134 3677 7146 3729
rect 7198 3677 7204 3729
rect 7012 3664 7204 3677
rect 7012 2972 7018 3664
rect 7198 2972 7204 3664
rect 7012 2969 7019 2972
rect 7053 2969 7091 2972
rect 7125 2969 7163 2972
rect 7197 2969 7204 2972
rect 7012 2930 7204 2969
rect 7012 2896 7019 2930
rect 7053 2896 7091 2930
rect 7125 2896 7163 2930
rect 7197 2896 7204 2930
rect 7012 2857 7204 2896
rect 7012 2823 7019 2857
rect 7053 2823 7091 2857
rect 7125 2823 7163 2857
rect 7197 2823 7204 2857
rect 7012 2784 7204 2823
rect 7012 2750 7019 2784
rect 7053 2750 7091 2784
rect 7125 2750 7163 2784
rect 7197 2750 7204 2784
rect 7012 2711 7204 2750
rect 7012 2677 7019 2711
rect 7053 2677 7091 2711
rect 7125 2677 7163 2711
rect 7197 2677 7204 2711
rect 7012 2638 7204 2677
rect 7012 2604 7019 2638
rect 7053 2604 7091 2638
rect 7125 2604 7163 2638
rect 7197 2604 7204 2638
rect 7012 2565 7204 2604
rect 7012 2531 7019 2565
rect 7053 2531 7091 2565
rect 7125 2531 7163 2565
rect 7197 2531 7204 2565
rect 7012 2492 7204 2531
rect 7012 2458 7019 2492
rect 7053 2458 7091 2492
rect 7125 2458 7163 2492
rect 7197 2458 7204 2492
rect 7012 2419 7204 2458
rect 7012 2385 7019 2419
rect 7053 2385 7091 2419
rect 7125 2385 7163 2419
rect 7197 2385 7204 2419
rect 7012 2346 7204 2385
rect 7012 2312 7019 2346
rect 7053 2312 7091 2346
rect 7125 2312 7163 2346
rect 7197 2312 7204 2346
rect 7012 2273 7204 2312
rect 7012 2239 7019 2273
rect 7053 2239 7091 2273
rect 7125 2239 7163 2273
rect 7197 2239 7204 2273
rect 7012 2200 7204 2239
rect 7012 2166 7019 2200
rect 7053 2166 7091 2200
rect 7125 2166 7163 2200
rect 7197 2166 7204 2200
rect 7012 2126 7204 2166
rect 7012 2092 7019 2126
rect 7053 2092 7091 2126
rect 7125 2092 7163 2126
rect 7197 2092 7204 2126
rect 7012 2052 7204 2092
rect 7012 2018 7019 2052
rect 7053 2018 7091 2052
rect 7125 2018 7163 2052
rect 7197 2018 7204 2052
rect 7012 1978 7204 2018
rect 7012 1944 7019 1978
rect 7053 1944 7091 1978
rect 7125 1944 7163 1978
rect 7197 1944 7204 1978
rect 7012 1904 7204 1944
rect 7012 1870 7019 1904
rect 7053 1870 7091 1904
rect 7125 1870 7163 1904
rect 7197 1870 7204 1904
rect 7012 1830 7204 1870
rect 7012 1796 7019 1830
rect 7053 1796 7091 1830
rect 7125 1796 7163 1830
rect 7197 1796 7204 1830
rect 7012 1756 7204 1796
rect 7012 1722 7019 1756
rect 7053 1722 7091 1756
rect 7125 1722 7163 1756
rect 7197 1722 7204 1756
rect 7012 1682 7204 1722
rect 7012 1648 7019 1682
rect 7053 1648 7091 1682
rect 7125 1648 7163 1682
rect 7197 1648 7204 1682
rect 7012 1608 7204 1648
rect 7012 1574 7019 1608
rect 7053 1574 7091 1608
rect 7125 1574 7163 1608
rect 7197 1574 7204 1608
rect 7012 1562 7204 1574
rect 7508 4118 7700 4130
rect 7508 4092 7587 4118
rect 7621 4092 7700 4118
rect 7508 3194 7515 4092
rect 7693 3194 7700 4092
rect 7508 3182 7700 3194
rect 7508 3148 7587 3182
rect 7621 3148 7700 3182
rect 7508 3108 7700 3148
rect 7508 3074 7515 3108
rect 7549 3074 7587 3108
rect 7621 3074 7659 3108
rect 7693 3074 7700 3108
rect 7508 3028 7700 3074
rect 7508 2994 7515 3028
rect 7549 2994 7587 3028
rect 7621 2994 7659 3028
rect 7693 2994 7700 3028
rect 7508 2948 7700 2994
rect 7508 2914 7515 2948
rect 7549 2914 7587 2948
rect 7621 2914 7659 2948
rect 7693 2914 7700 2948
rect 7508 2868 7700 2914
rect 7508 2834 7515 2868
rect 7549 2834 7587 2868
rect 7621 2834 7659 2868
rect 7693 2834 7700 2868
rect 7508 2788 7700 2834
rect 7508 2754 7515 2788
rect 7549 2754 7587 2788
rect 7621 2754 7659 2788
rect 7693 2754 7700 2788
rect 7508 2708 7700 2754
rect 7508 2674 7515 2708
rect 7549 2674 7587 2708
rect 7621 2674 7659 2708
rect 7693 2674 7700 2708
rect 7508 2657 7700 2674
rect 7508 2605 7514 2657
rect 7566 2605 7578 2657
rect 7630 2605 7642 2657
rect 7694 2605 7700 2657
rect 7508 2594 7515 2605
rect 7549 2594 7587 2605
rect 7621 2594 7659 2605
rect 7693 2594 7700 2605
rect 7508 2592 7700 2594
rect 7508 2540 7514 2592
rect 7566 2540 7578 2592
rect 7630 2540 7642 2592
rect 7694 2540 7700 2592
rect 7508 2527 7587 2540
rect 7621 2527 7700 2540
rect 7508 2475 7514 2527
rect 7566 2518 7578 2527
rect 7630 2518 7642 2527
rect 7694 2475 7700 2527
rect 7508 2462 7515 2475
rect 7693 2462 7700 2475
rect 7508 2410 7514 2462
rect 7694 2410 7700 2462
rect 7508 2397 7515 2410
rect 7693 2397 7700 2410
rect 7508 2345 7514 2397
rect 7694 2345 7700 2397
rect 7508 2332 7515 2345
rect 7693 2332 7700 2345
rect 7508 2280 7514 2332
rect 7694 2280 7700 2332
rect 7508 2267 7515 2280
rect 7693 2267 7700 2280
rect 7508 2215 7514 2267
rect 7694 2215 7700 2267
rect 7508 2202 7515 2215
rect 7693 2202 7700 2215
rect 7508 2150 7514 2202
rect 7694 2150 7700 2202
rect 7508 2137 7515 2150
rect 7693 2137 7700 2150
rect 7508 2085 7514 2137
rect 7694 2085 7700 2137
rect 7508 2072 7515 2085
rect 7693 2072 7700 2085
rect 7508 2020 7514 2072
rect 7694 2020 7700 2072
rect 7508 2007 7515 2020
rect 7693 2007 7700 2020
rect 7508 1955 7514 2007
rect 7694 1955 7700 2007
rect 7508 1942 7515 1955
rect 7693 1942 7700 1955
rect 7508 1890 7514 1942
rect 7694 1890 7700 1942
rect 7508 1877 7515 1890
rect 7693 1877 7700 1890
rect 7508 1825 7514 1877
rect 7694 1825 7700 1877
rect 7508 1812 7515 1825
rect 7693 1812 7700 1825
rect 7508 1568 7514 1812
rect 7694 1568 7700 1812
rect 7508 1562 7700 1568
rect 8004 4119 8196 4125
rect 8004 4067 8010 4119
rect 8062 4067 8074 4119
rect 8126 4067 8138 4119
rect 8190 4067 8196 4119
rect 8004 4064 8011 4067
rect 8045 4064 8083 4067
rect 8117 4064 8155 4067
rect 8189 4064 8196 4067
rect 8004 4054 8196 4064
rect 8004 4002 8010 4054
rect 8062 4002 8074 4054
rect 8126 4002 8138 4054
rect 8190 4002 8196 4054
rect 8004 3991 8011 4002
rect 8045 3991 8083 4002
rect 8117 3991 8155 4002
rect 8189 3991 8196 4002
rect 8004 3989 8196 3991
rect 8004 3937 8010 3989
rect 8062 3937 8074 3989
rect 8126 3937 8138 3989
rect 8190 3937 8196 3989
rect 8004 3924 8011 3937
rect 8045 3924 8083 3937
rect 8117 3924 8155 3937
rect 8189 3924 8196 3937
rect 8004 3872 8010 3924
rect 8062 3872 8074 3924
rect 8126 3872 8138 3924
rect 8190 3872 8196 3924
rect 8004 3859 8011 3872
rect 8045 3859 8083 3872
rect 8117 3859 8155 3872
rect 8189 3859 8196 3872
rect 8004 3807 8010 3859
rect 8062 3807 8074 3859
rect 8126 3807 8138 3859
rect 8190 3807 8196 3859
rect 8004 3806 8196 3807
rect 8004 3794 8011 3806
rect 8045 3794 8083 3806
rect 8117 3794 8155 3806
rect 8189 3794 8196 3806
rect 8004 3742 8010 3794
rect 8062 3742 8074 3794
rect 8126 3742 8138 3794
rect 8190 3742 8196 3794
rect 8004 3733 8196 3742
rect 8004 3729 8011 3733
rect 8045 3729 8083 3733
rect 8117 3729 8155 3733
rect 8189 3729 8196 3733
rect 8004 3677 8010 3729
rect 8062 3677 8074 3729
rect 8126 3677 8138 3729
rect 8190 3677 8196 3729
rect 8004 3664 8196 3677
rect 8004 2972 8010 3664
rect 8190 2972 8196 3664
rect 8004 2969 8011 2972
rect 8045 2969 8083 2972
rect 8117 2969 8155 2972
rect 8189 2969 8196 2972
rect 8004 2930 8196 2969
rect 8004 2896 8011 2930
rect 8045 2896 8083 2930
rect 8117 2896 8155 2930
rect 8189 2896 8196 2930
rect 8004 2857 8196 2896
rect 8004 2823 8011 2857
rect 8045 2823 8083 2857
rect 8117 2823 8155 2857
rect 8189 2823 8196 2857
rect 8004 2784 8196 2823
rect 8004 2750 8011 2784
rect 8045 2750 8083 2784
rect 8117 2750 8155 2784
rect 8189 2750 8196 2784
rect 8004 2711 8196 2750
rect 8004 2677 8011 2711
rect 8045 2677 8083 2711
rect 8117 2677 8155 2711
rect 8189 2677 8196 2711
rect 8004 2638 8196 2677
rect 8004 2604 8011 2638
rect 8045 2604 8083 2638
rect 8117 2604 8155 2638
rect 8189 2604 8196 2638
rect 8004 2565 8196 2604
rect 8004 2531 8011 2565
rect 8045 2531 8083 2565
rect 8117 2531 8155 2565
rect 8189 2531 8196 2565
rect 8004 2492 8196 2531
rect 8004 2458 8011 2492
rect 8045 2458 8083 2492
rect 8117 2458 8155 2492
rect 8189 2458 8196 2492
rect 8004 2419 8196 2458
rect 8004 2385 8011 2419
rect 8045 2385 8083 2419
rect 8117 2385 8155 2419
rect 8189 2385 8196 2419
rect 8004 2346 8196 2385
rect 8004 2312 8011 2346
rect 8045 2312 8083 2346
rect 8117 2312 8155 2346
rect 8189 2312 8196 2346
rect 8004 2273 8196 2312
rect 8004 2239 8011 2273
rect 8045 2239 8083 2273
rect 8117 2239 8155 2273
rect 8189 2239 8196 2273
rect 8004 2200 8196 2239
rect 8004 2166 8011 2200
rect 8045 2166 8083 2200
rect 8117 2166 8155 2200
rect 8189 2166 8196 2200
rect 8004 2126 8196 2166
rect 8004 2092 8011 2126
rect 8045 2092 8083 2126
rect 8117 2092 8155 2126
rect 8189 2092 8196 2126
rect 8004 2052 8196 2092
rect 8004 2018 8011 2052
rect 8045 2018 8083 2052
rect 8117 2018 8155 2052
rect 8189 2018 8196 2052
rect 8004 1978 8196 2018
rect 8004 1944 8011 1978
rect 8045 1944 8083 1978
rect 8117 1944 8155 1978
rect 8189 1944 8196 1978
rect 8004 1904 8196 1944
rect 8004 1870 8011 1904
rect 8045 1870 8083 1904
rect 8117 1870 8155 1904
rect 8189 1870 8196 1904
rect 8004 1830 8196 1870
rect 8004 1796 8011 1830
rect 8045 1796 8083 1830
rect 8117 1796 8155 1830
rect 8189 1796 8196 1830
rect 8004 1756 8196 1796
rect 8004 1722 8011 1756
rect 8045 1722 8083 1756
rect 8117 1722 8155 1756
rect 8189 1722 8196 1756
rect 8004 1682 8196 1722
rect 8004 1648 8011 1682
rect 8045 1648 8083 1682
rect 8117 1648 8155 1682
rect 8189 1648 8196 1682
rect 8004 1608 8196 1648
rect 8004 1574 8011 1608
rect 8045 1574 8083 1608
rect 8117 1574 8155 1608
rect 8189 1574 8196 1608
rect 8004 1562 8196 1574
rect 8500 4118 8692 4130
rect 8500 4092 8579 4118
rect 8613 4092 8692 4118
rect 8500 3194 8507 4092
rect 8685 3194 8692 4092
rect 8500 3182 8692 3194
rect 8500 3148 8579 3182
rect 8613 3148 8692 3182
rect 8500 3108 8692 3148
rect 8500 3074 8507 3108
rect 8541 3074 8579 3108
rect 8613 3074 8651 3108
rect 8685 3074 8692 3108
rect 8500 3028 8692 3074
rect 8500 2994 8507 3028
rect 8541 2994 8579 3028
rect 8613 2994 8651 3028
rect 8685 2994 8692 3028
rect 8500 2948 8692 2994
rect 8500 2914 8507 2948
rect 8541 2914 8579 2948
rect 8613 2914 8651 2948
rect 8685 2914 8692 2948
rect 8500 2868 8692 2914
rect 8500 2834 8507 2868
rect 8541 2834 8579 2868
rect 8613 2834 8651 2868
rect 8685 2834 8692 2868
rect 8500 2788 8692 2834
rect 8500 2754 8507 2788
rect 8541 2754 8579 2788
rect 8613 2754 8651 2788
rect 8685 2754 8692 2788
rect 8500 2708 8692 2754
rect 8500 2674 8507 2708
rect 8541 2674 8579 2708
rect 8613 2674 8651 2708
rect 8685 2674 8692 2708
rect 8500 2657 8692 2674
rect 8500 2605 8506 2657
rect 8558 2605 8570 2657
rect 8622 2605 8634 2657
rect 8686 2605 8692 2657
rect 8500 2594 8507 2605
rect 8541 2594 8579 2605
rect 8613 2594 8651 2605
rect 8685 2594 8692 2605
rect 8500 2592 8692 2594
rect 8500 2540 8506 2592
rect 8558 2540 8570 2592
rect 8622 2540 8634 2592
rect 8686 2540 8692 2592
rect 8500 2527 8579 2540
rect 8613 2527 8692 2540
rect 8500 2475 8506 2527
rect 8558 2518 8570 2527
rect 8622 2518 8634 2527
rect 8686 2475 8692 2527
rect 8500 2462 8507 2475
rect 8685 2462 8692 2475
rect 8500 2410 8506 2462
rect 8686 2410 8692 2462
rect 8500 2397 8507 2410
rect 8685 2397 8692 2410
rect 8500 2345 8506 2397
rect 8686 2345 8692 2397
rect 8500 2332 8507 2345
rect 8685 2332 8692 2345
rect 8500 2280 8506 2332
rect 8686 2280 8692 2332
rect 8500 2267 8507 2280
rect 8685 2267 8692 2280
rect 8500 2215 8506 2267
rect 8686 2215 8692 2267
rect 8500 2202 8507 2215
rect 8685 2202 8692 2215
rect 8500 2150 8506 2202
rect 8686 2150 8692 2202
rect 8500 2137 8507 2150
rect 8685 2137 8692 2150
rect 8500 2085 8506 2137
rect 8686 2085 8692 2137
rect 8500 2072 8507 2085
rect 8685 2072 8692 2085
rect 8500 2020 8506 2072
rect 8686 2020 8692 2072
rect 8500 2007 8507 2020
rect 8685 2007 8692 2020
rect 8500 1955 8506 2007
rect 8686 1955 8692 2007
rect 8500 1942 8507 1955
rect 8685 1942 8692 1955
rect 8500 1890 8506 1942
rect 8686 1890 8692 1942
rect 8500 1877 8507 1890
rect 8685 1877 8692 1890
rect 8500 1825 8506 1877
rect 8686 1825 8692 1877
rect 8500 1812 8507 1825
rect 8685 1812 8692 1825
rect 8500 1568 8506 1812
rect 8686 1568 8692 1812
rect 8500 1562 8692 1568
rect 8996 4119 9188 4125
rect 8996 4067 9002 4119
rect 9054 4067 9066 4119
rect 9118 4067 9130 4119
rect 9182 4067 9188 4119
rect 8996 4064 9003 4067
rect 9037 4064 9075 4067
rect 9109 4064 9147 4067
rect 9181 4064 9188 4067
rect 8996 4054 9188 4064
rect 8996 4002 9002 4054
rect 9054 4002 9066 4054
rect 9118 4002 9130 4054
rect 9182 4002 9188 4054
rect 8996 3991 9003 4002
rect 9037 3991 9075 4002
rect 9109 3991 9147 4002
rect 9181 3991 9188 4002
rect 8996 3989 9188 3991
rect 8996 3937 9002 3989
rect 9054 3937 9066 3989
rect 9118 3937 9130 3989
rect 9182 3937 9188 3989
rect 8996 3924 9003 3937
rect 9037 3924 9075 3937
rect 9109 3924 9147 3937
rect 9181 3924 9188 3937
rect 8996 3872 9002 3924
rect 9054 3872 9066 3924
rect 9118 3872 9130 3924
rect 9182 3872 9188 3924
rect 8996 3859 9003 3872
rect 9037 3859 9075 3872
rect 9109 3859 9147 3872
rect 9181 3859 9188 3872
rect 8996 3807 9002 3859
rect 9054 3807 9066 3859
rect 9118 3807 9130 3859
rect 9182 3807 9188 3859
rect 8996 3806 9188 3807
rect 8996 3794 9003 3806
rect 9037 3794 9075 3806
rect 9109 3794 9147 3806
rect 9181 3794 9188 3806
rect 8996 3742 9002 3794
rect 9054 3742 9066 3794
rect 9118 3742 9130 3794
rect 9182 3742 9188 3794
rect 8996 3733 9188 3742
rect 8996 3729 9003 3733
rect 9037 3729 9075 3733
rect 9109 3729 9147 3733
rect 9181 3729 9188 3733
rect 8996 3677 9002 3729
rect 9054 3677 9066 3729
rect 9118 3677 9130 3729
rect 9182 3677 9188 3729
rect 8996 3664 9188 3677
rect 8996 2972 9002 3664
rect 9182 2972 9188 3664
rect 8996 2969 9003 2972
rect 9037 2969 9075 2972
rect 9109 2969 9147 2972
rect 9181 2969 9188 2972
rect 8996 2930 9188 2969
rect 8996 2896 9003 2930
rect 9037 2896 9075 2930
rect 9109 2896 9147 2930
rect 9181 2896 9188 2930
rect 8996 2857 9188 2896
rect 8996 2823 9003 2857
rect 9037 2823 9075 2857
rect 9109 2823 9147 2857
rect 9181 2823 9188 2857
rect 8996 2784 9188 2823
rect 8996 2750 9003 2784
rect 9037 2750 9075 2784
rect 9109 2750 9147 2784
rect 9181 2750 9188 2784
rect 8996 2711 9188 2750
rect 8996 2677 9003 2711
rect 9037 2677 9075 2711
rect 9109 2677 9147 2711
rect 9181 2677 9188 2711
rect 8996 2638 9188 2677
rect 8996 2604 9003 2638
rect 9037 2604 9075 2638
rect 9109 2604 9147 2638
rect 9181 2604 9188 2638
rect 8996 2565 9188 2604
rect 8996 2531 9003 2565
rect 9037 2531 9075 2565
rect 9109 2531 9147 2565
rect 9181 2531 9188 2565
rect 8996 2492 9188 2531
rect 8996 2458 9003 2492
rect 9037 2458 9075 2492
rect 9109 2458 9147 2492
rect 9181 2458 9188 2492
rect 8996 2419 9188 2458
rect 8996 2385 9003 2419
rect 9037 2385 9075 2419
rect 9109 2385 9147 2419
rect 9181 2385 9188 2419
rect 8996 2346 9188 2385
rect 8996 2312 9003 2346
rect 9037 2312 9075 2346
rect 9109 2312 9147 2346
rect 9181 2312 9188 2346
rect 8996 2273 9188 2312
rect 8996 2239 9003 2273
rect 9037 2239 9075 2273
rect 9109 2239 9147 2273
rect 9181 2239 9188 2273
rect 8996 2200 9188 2239
rect 8996 2166 9003 2200
rect 9037 2166 9075 2200
rect 9109 2166 9147 2200
rect 9181 2166 9188 2200
rect 8996 2126 9188 2166
rect 8996 2092 9003 2126
rect 9037 2092 9075 2126
rect 9109 2092 9147 2126
rect 9181 2092 9188 2126
rect 8996 2052 9188 2092
rect 8996 2018 9003 2052
rect 9037 2018 9075 2052
rect 9109 2018 9147 2052
rect 9181 2018 9188 2052
rect 8996 1978 9188 2018
rect 8996 1944 9003 1978
rect 9037 1944 9075 1978
rect 9109 1944 9147 1978
rect 9181 1944 9188 1978
rect 8996 1904 9188 1944
rect 8996 1870 9003 1904
rect 9037 1870 9075 1904
rect 9109 1870 9147 1904
rect 9181 1870 9188 1904
rect 8996 1830 9188 1870
rect 8996 1796 9003 1830
rect 9037 1796 9075 1830
rect 9109 1796 9147 1830
rect 9181 1796 9188 1830
rect 8996 1756 9188 1796
rect 8996 1722 9003 1756
rect 9037 1722 9075 1756
rect 9109 1722 9147 1756
rect 9181 1722 9188 1756
rect 8996 1682 9188 1722
rect 8996 1648 9003 1682
rect 9037 1648 9075 1682
rect 9109 1648 9147 1682
rect 9181 1648 9188 1682
rect 8996 1608 9188 1648
rect 8996 1574 9003 1608
rect 9037 1574 9075 1608
rect 9109 1574 9147 1608
rect 9181 1574 9188 1608
rect 8996 1562 9188 1574
rect 9492 4118 9684 4130
rect 9492 4092 9571 4118
rect 9605 4092 9684 4118
rect 9492 3194 9499 4092
rect 9677 3194 9684 4092
rect 9492 3182 9684 3194
rect 9492 3148 9571 3182
rect 9605 3148 9684 3182
rect 9492 3108 9684 3148
rect 9492 3074 9499 3108
rect 9533 3074 9571 3108
rect 9605 3074 9643 3108
rect 9677 3074 9684 3108
rect 9492 3028 9684 3074
rect 9492 2994 9499 3028
rect 9533 2994 9571 3028
rect 9605 2994 9643 3028
rect 9677 2994 9684 3028
rect 9492 2948 9684 2994
rect 9492 2914 9499 2948
rect 9533 2914 9571 2948
rect 9605 2914 9643 2948
rect 9677 2914 9684 2948
rect 9492 2868 9684 2914
rect 9492 2834 9499 2868
rect 9533 2834 9571 2868
rect 9605 2834 9643 2868
rect 9677 2834 9684 2868
rect 9492 2788 9684 2834
rect 9492 2754 9499 2788
rect 9533 2754 9571 2788
rect 9605 2754 9643 2788
rect 9677 2754 9684 2788
rect 9492 2708 9684 2754
rect 9492 2674 9499 2708
rect 9533 2674 9571 2708
rect 9605 2674 9643 2708
rect 9677 2674 9684 2708
rect 9492 2657 9684 2674
rect 9492 2605 9498 2657
rect 9550 2605 9562 2657
rect 9614 2605 9626 2657
rect 9678 2605 9684 2657
rect 9492 2594 9499 2605
rect 9533 2594 9571 2605
rect 9605 2594 9643 2605
rect 9677 2594 9684 2605
rect 9492 2592 9684 2594
rect 9492 2540 9498 2592
rect 9550 2540 9562 2592
rect 9614 2540 9626 2592
rect 9678 2540 9684 2592
rect 9492 2527 9571 2540
rect 9605 2527 9684 2540
rect 9492 2475 9498 2527
rect 9550 2518 9562 2527
rect 9614 2518 9626 2527
rect 9678 2475 9684 2527
rect 9492 2462 9499 2475
rect 9677 2462 9684 2475
rect 9492 2410 9498 2462
rect 9678 2410 9684 2462
rect 9492 2397 9499 2410
rect 9677 2397 9684 2410
rect 9492 2345 9498 2397
rect 9678 2345 9684 2397
rect 9492 2332 9499 2345
rect 9677 2332 9684 2345
rect 9492 2280 9498 2332
rect 9678 2280 9684 2332
rect 9492 2267 9499 2280
rect 9677 2267 9684 2280
rect 9492 2215 9498 2267
rect 9678 2215 9684 2267
rect 9492 2202 9499 2215
rect 9677 2202 9684 2215
rect 9492 2150 9498 2202
rect 9678 2150 9684 2202
rect 9492 2137 9499 2150
rect 9677 2137 9684 2150
rect 9492 2085 9498 2137
rect 9678 2085 9684 2137
rect 9492 2072 9499 2085
rect 9677 2072 9684 2085
rect 9492 2020 9498 2072
rect 9678 2020 9684 2072
rect 9492 2007 9499 2020
rect 9677 2007 9684 2020
rect 9492 1955 9498 2007
rect 9678 1955 9684 2007
rect 9492 1942 9499 1955
rect 9677 1942 9684 1955
rect 9492 1890 9498 1942
rect 9678 1890 9684 1942
rect 9492 1877 9499 1890
rect 9677 1877 9684 1890
rect 9492 1825 9498 1877
rect 9678 1825 9684 1877
rect 9492 1812 9499 1825
rect 9677 1812 9684 1825
rect 9492 1568 9498 1812
rect 9678 1568 9684 1812
rect 9492 1562 9684 1568
rect 9988 4119 10180 4125
rect 9988 4067 9994 4119
rect 10046 4067 10058 4119
rect 10110 4067 10122 4119
rect 10174 4067 10180 4119
rect 9988 4064 9995 4067
rect 10029 4064 10067 4067
rect 10101 4064 10139 4067
rect 10173 4064 10180 4067
rect 9988 4054 10180 4064
rect 9988 4002 9994 4054
rect 10046 4002 10058 4054
rect 10110 4002 10122 4054
rect 10174 4002 10180 4054
rect 9988 3991 9995 4002
rect 10029 3991 10067 4002
rect 10101 3991 10139 4002
rect 10173 3991 10180 4002
rect 9988 3989 10180 3991
rect 9988 3937 9994 3989
rect 10046 3937 10058 3989
rect 10110 3937 10122 3989
rect 10174 3937 10180 3989
rect 9988 3924 9995 3937
rect 10029 3924 10067 3937
rect 10101 3924 10139 3937
rect 10173 3924 10180 3937
rect 9988 3872 9994 3924
rect 10046 3872 10058 3924
rect 10110 3872 10122 3924
rect 10174 3872 10180 3924
rect 9988 3859 9995 3872
rect 10029 3859 10067 3872
rect 10101 3859 10139 3872
rect 10173 3859 10180 3872
rect 9988 3807 9994 3859
rect 10046 3807 10058 3859
rect 10110 3807 10122 3859
rect 10174 3807 10180 3859
rect 9988 3806 10180 3807
rect 9988 3794 9995 3806
rect 10029 3794 10067 3806
rect 10101 3794 10139 3806
rect 10173 3794 10180 3806
rect 9988 3742 9994 3794
rect 10046 3742 10058 3794
rect 10110 3742 10122 3794
rect 10174 3742 10180 3794
rect 9988 3733 10180 3742
rect 9988 3729 9995 3733
rect 10029 3729 10067 3733
rect 10101 3729 10139 3733
rect 10173 3729 10180 3733
rect 9988 3677 9994 3729
rect 10046 3677 10058 3729
rect 10110 3677 10122 3729
rect 10174 3677 10180 3729
rect 9988 3664 10180 3677
rect 9988 2972 9994 3664
rect 10174 2972 10180 3664
rect 9988 2969 9995 2972
rect 10029 2969 10067 2972
rect 10101 2969 10139 2972
rect 10173 2969 10180 2972
rect 9988 2930 10180 2969
rect 9988 2896 9995 2930
rect 10029 2896 10067 2930
rect 10101 2896 10139 2930
rect 10173 2896 10180 2930
rect 9988 2857 10180 2896
rect 9988 2823 9995 2857
rect 10029 2823 10067 2857
rect 10101 2823 10139 2857
rect 10173 2823 10180 2857
rect 9988 2784 10180 2823
rect 9988 2750 9995 2784
rect 10029 2750 10067 2784
rect 10101 2750 10139 2784
rect 10173 2750 10180 2784
rect 9988 2711 10180 2750
rect 9988 2677 9995 2711
rect 10029 2677 10067 2711
rect 10101 2677 10139 2711
rect 10173 2677 10180 2711
rect 9988 2638 10180 2677
rect 9988 2604 9995 2638
rect 10029 2604 10067 2638
rect 10101 2604 10139 2638
rect 10173 2604 10180 2638
rect 9988 2565 10180 2604
rect 9988 2531 9995 2565
rect 10029 2531 10067 2565
rect 10101 2531 10139 2565
rect 10173 2531 10180 2565
rect 9988 2492 10180 2531
rect 9988 2458 9995 2492
rect 10029 2458 10067 2492
rect 10101 2458 10139 2492
rect 10173 2458 10180 2492
rect 9988 2419 10180 2458
rect 9988 2385 9995 2419
rect 10029 2385 10067 2419
rect 10101 2385 10139 2419
rect 10173 2385 10180 2419
rect 9988 2346 10180 2385
rect 9988 2312 9995 2346
rect 10029 2312 10067 2346
rect 10101 2312 10139 2346
rect 10173 2312 10180 2346
rect 9988 2273 10180 2312
rect 9988 2239 9995 2273
rect 10029 2239 10067 2273
rect 10101 2239 10139 2273
rect 10173 2239 10180 2273
rect 9988 2200 10180 2239
rect 9988 2166 9995 2200
rect 10029 2166 10067 2200
rect 10101 2166 10139 2200
rect 10173 2166 10180 2200
rect 9988 2126 10180 2166
rect 9988 2092 9995 2126
rect 10029 2092 10067 2126
rect 10101 2092 10139 2126
rect 10173 2092 10180 2126
rect 9988 2052 10180 2092
rect 9988 2018 9995 2052
rect 10029 2018 10067 2052
rect 10101 2018 10139 2052
rect 10173 2018 10180 2052
rect 9988 1978 10180 2018
rect 9988 1944 9995 1978
rect 10029 1944 10067 1978
rect 10101 1944 10139 1978
rect 10173 1944 10180 1978
rect 9988 1904 10180 1944
rect 9988 1870 9995 1904
rect 10029 1870 10067 1904
rect 10101 1870 10139 1904
rect 10173 1870 10180 1904
rect 9988 1830 10180 1870
rect 9988 1796 9995 1830
rect 10029 1796 10067 1830
rect 10101 1796 10139 1830
rect 10173 1796 10180 1830
rect 9988 1756 10180 1796
rect 9988 1722 9995 1756
rect 10029 1722 10067 1756
rect 10101 1722 10139 1756
rect 10173 1722 10180 1756
rect 9988 1682 10180 1722
rect 9988 1648 9995 1682
rect 10029 1648 10067 1682
rect 10101 1648 10139 1682
rect 10173 1648 10180 1682
rect 9988 1608 10180 1648
rect 9988 1574 9995 1608
rect 10029 1574 10067 1608
rect 10101 1574 10139 1608
rect 10173 1574 10180 1608
rect 9988 1562 10180 1574
rect 10484 4118 10676 4130
rect 10484 4092 10563 4118
rect 10597 4092 10676 4118
rect 10484 3194 10491 4092
rect 10669 3194 10676 4092
rect 10484 3182 10676 3194
rect 10484 3148 10563 3182
rect 10597 3148 10676 3182
rect 10484 3108 10676 3148
rect 10484 3074 10491 3108
rect 10525 3074 10563 3108
rect 10597 3074 10635 3108
rect 10669 3074 10676 3108
rect 10484 3028 10676 3074
rect 10484 2994 10491 3028
rect 10525 2994 10563 3028
rect 10597 2994 10635 3028
rect 10669 2994 10676 3028
rect 10484 2948 10676 2994
rect 10484 2914 10491 2948
rect 10525 2914 10563 2948
rect 10597 2914 10635 2948
rect 10669 2914 10676 2948
rect 10484 2868 10676 2914
rect 10484 2834 10491 2868
rect 10525 2834 10563 2868
rect 10597 2834 10635 2868
rect 10669 2834 10676 2868
rect 10484 2788 10676 2834
rect 10484 2754 10491 2788
rect 10525 2754 10563 2788
rect 10597 2754 10635 2788
rect 10669 2754 10676 2788
rect 10484 2708 10676 2754
rect 10484 2674 10491 2708
rect 10525 2674 10563 2708
rect 10597 2674 10635 2708
rect 10669 2674 10676 2708
rect 10484 2657 10676 2674
rect 10484 2605 10490 2657
rect 10542 2605 10554 2657
rect 10606 2605 10618 2657
rect 10670 2605 10676 2657
rect 10484 2594 10491 2605
rect 10525 2594 10563 2605
rect 10597 2594 10635 2605
rect 10669 2594 10676 2605
rect 10484 2592 10676 2594
rect 10484 2540 10490 2592
rect 10542 2540 10554 2592
rect 10606 2540 10618 2592
rect 10670 2540 10676 2592
rect 10484 2527 10563 2540
rect 10597 2527 10676 2540
rect 10484 2475 10490 2527
rect 10542 2518 10554 2527
rect 10606 2518 10618 2527
rect 10670 2475 10676 2527
rect 10484 2462 10491 2475
rect 10669 2462 10676 2475
rect 10484 2410 10490 2462
rect 10670 2410 10676 2462
rect 10484 2397 10491 2410
rect 10669 2397 10676 2410
rect 10484 2345 10490 2397
rect 10670 2345 10676 2397
rect 10484 2332 10491 2345
rect 10669 2332 10676 2345
rect 10484 2280 10490 2332
rect 10670 2280 10676 2332
rect 10484 2267 10491 2280
rect 10669 2267 10676 2280
rect 10484 2215 10490 2267
rect 10670 2215 10676 2267
rect 10484 2202 10491 2215
rect 10669 2202 10676 2215
rect 10484 2150 10490 2202
rect 10670 2150 10676 2202
rect 10484 2137 10491 2150
rect 10669 2137 10676 2150
rect 10484 2085 10490 2137
rect 10670 2085 10676 2137
rect 10484 2072 10491 2085
rect 10669 2072 10676 2085
rect 10484 2020 10490 2072
rect 10670 2020 10676 2072
rect 10484 2007 10491 2020
rect 10669 2007 10676 2020
rect 10484 1955 10490 2007
rect 10670 1955 10676 2007
rect 10484 1942 10491 1955
rect 10669 1942 10676 1955
rect 10484 1890 10490 1942
rect 10670 1890 10676 1942
rect 10484 1877 10491 1890
rect 10669 1877 10676 1890
rect 10484 1825 10490 1877
rect 10670 1825 10676 1877
rect 10484 1812 10491 1825
rect 10669 1812 10676 1825
rect 10484 1568 10490 1812
rect 10670 1568 10676 1812
rect 10484 1562 10676 1568
rect 10980 4119 11172 4125
rect 10980 4067 10986 4119
rect 11038 4067 11050 4119
rect 11102 4067 11114 4119
rect 11166 4067 11172 4119
rect 10980 4064 10987 4067
rect 11021 4064 11059 4067
rect 11093 4064 11131 4067
rect 11165 4064 11172 4067
rect 10980 4054 11172 4064
rect 10980 4002 10986 4054
rect 11038 4002 11050 4054
rect 11102 4002 11114 4054
rect 11166 4002 11172 4054
rect 10980 3991 10987 4002
rect 11021 3991 11059 4002
rect 11093 3991 11131 4002
rect 11165 3991 11172 4002
rect 10980 3989 11172 3991
rect 10980 3937 10986 3989
rect 11038 3937 11050 3989
rect 11102 3937 11114 3989
rect 11166 3937 11172 3989
rect 10980 3924 10987 3937
rect 11021 3924 11059 3937
rect 11093 3924 11131 3937
rect 11165 3924 11172 3937
rect 10980 3872 10986 3924
rect 11038 3872 11050 3924
rect 11102 3872 11114 3924
rect 11166 3872 11172 3924
rect 10980 3859 10987 3872
rect 11021 3859 11059 3872
rect 11093 3859 11131 3872
rect 11165 3859 11172 3872
rect 10980 3807 10986 3859
rect 11038 3807 11050 3859
rect 11102 3807 11114 3859
rect 11166 3807 11172 3859
rect 10980 3806 11172 3807
rect 10980 3794 10987 3806
rect 11021 3794 11059 3806
rect 11093 3794 11131 3806
rect 11165 3794 11172 3806
rect 10980 3742 10986 3794
rect 11038 3742 11050 3794
rect 11102 3742 11114 3794
rect 11166 3742 11172 3794
rect 10980 3733 11172 3742
rect 10980 3729 10987 3733
rect 11021 3729 11059 3733
rect 11093 3729 11131 3733
rect 11165 3729 11172 3733
rect 10980 3677 10986 3729
rect 11038 3677 11050 3729
rect 11102 3677 11114 3729
rect 11166 3677 11172 3729
rect 10980 3664 11172 3677
rect 10980 2972 10986 3664
rect 11166 2972 11172 3664
rect 10980 2969 10987 2972
rect 11021 2969 11059 2972
rect 11093 2969 11131 2972
rect 11165 2969 11172 2972
rect 10980 2930 11172 2969
rect 10980 2896 10987 2930
rect 11021 2896 11059 2930
rect 11093 2896 11131 2930
rect 11165 2896 11172 2930
rect 10980 2857 11172 2896
rect 10980 2823 10987 2857
rect 11021 2823 11059 2857
rect 11093 2823 11131 2857
rect 11165 2823 11172 2857
rect 10980 2784 11172 2823
rect 10980 2750 10987 2784
rect 11021 2750 11059 2784
rect 11093 2750 11131 2784
rect 11165 2750 11172 2784
rect 10980 2711 11172 2750
rect 10980 2677 10987 2711
rect 11021 2677 11059 2711
rect 11093 2677 11131 2711
rect 11165 2677 11172 2711
rect 10980 2638 11172 2677
rect 10980 2604 10987 2638
rect 11021 2604 11059 2638
rect 11093 2604 11131 2638
rect 11165 2604 11172 2638
rect 10980 2565 11172 2604
rect 10980 2531 10987 2565
rect 11021 2531 11059 2565
rect 11093 2531 11131 2565
rect 11165 2531 11172 2565
rect 10980 2492 11172 2531
rect 10980 2458 10987 2492
rect 11021 2458 11059 2492
rect 11093 2458 11131 2492
rect 11165 2458 11172 2492
rect 10980 2419 11172 2458
rect 10980 2385 10987 2419
rect 11021 2385 11059 2419
rect 11093 2385 11131 2419
rect 11165 2385 11172 2419
rect 10980 2346 11172 2385
rect 10980 2312 10987 2346
rect 11021 2312 11059 2346
rect 11093 2312 11131 2346
rect 11165 2312 11172 2346
rect 10980 2273 11172 2312
rect 10980 2239 10987 2273
rect 11021 2239 11059 2273
rect 11093 2239 11131 2273
rect 11165 2239 11172 2273
rect 10980 2200 11172 2239
rect 10980 2166 10987 2200
rect 11021 2166 11059 2200
rect 11093 2166 11131 2200
rect 11165 2166 11172 2200
rect 10980 2126 11172 2166
rect 10980 2092 10987 2126
rect 11021 2092 11059 2126
rect 11093 2092 11131 2126
rect 11165 2092 11172 2126
rect 10980 2052 11172 2092
rect 10980 2018 10987 2052
rect 11021 2018 11059 2052
rect 11093 2018 11131 2052
rect 11165 2018 11172 2052
rect 10980 1978 11172 2018
rect 10980 1944 10987 1978
rect 11021 1944 11059 1978
rect 11093 1944 11131 1978
rect 11165 1944 11172 1978
rect 10980 1904 11172 1944
rect 10980 1870 10987 1904
rect 11021 1870 11059 1904
rect 11093 1870 11131 1904
rect 11165 1870 11172 1904
rect 10980 1830 11172 1870
rect 10980 1796 10987 1830
rect 11021 1796 11059 1830
rect 11093 1796 11131 1830
rect 11165 1796 11172 1830
rect 10980 1756 11172 1796
rect 10980 1722 10987 1756
rect 11021 1722 11059 1756
rect 11093 1722 11131 1756
rect 11165 1722 11172 1756
rect 10980 1682 11172 1722
rect 10980 1648 10987 1682
rect 11021 1648 11059 1682
rect 11093 1648 11131 1682
rect 11165 1648 11172 1682
rect 10980 1608 11172 1648
rect 10980 1574 10987 1608
rect 11021 1574 11059 1608
rect 11093 1574 11131 1608
rect 11165 1574 11172 1608
rect 10980 1562 11172 1574
rect 11476 4118 11668 4130
rect 11476 4092 11555 4118
rect 11589 4092 11668 4118
rect 11476 3194 11483 4092
rect 11661 3194 11668 4092
rect 11476 3182 11668 3194
rect 11476 3148 11555 3182
rect 11589 3148 11668 3182
rect 11476 3108 11668 3148
rect 11476 3074 11483 3108
rect 11517 3074 11555 3108
rect 11589 3074 11627 3108
rect 11661 3074 11668 3108
rect 11476 3028 11668 3074
rect 11476 2994 11483 3028
rect 11517 2994 11555 3028
rect 11589 2994 11627 3028
rect 11661 2994 11668 3028
rect 11476 2948 11668 2994
rect 11476 2914 11483 2948
rect 11517 2914 11555 2948
rect 11589 2914 11627 2948
rect 11661 2914 11668 2948
rect 11476 2868 11668 2914
rect 11476 2834 11483 2868
rect 11517 2834 11555 2868
rect 11589 2834 11627 2868
rect 11661 2834 11668 2868
rect 11476 2788 11668 2834
rect 11476 2754 11483 2788
rect 11517 2754 11555 2788
rect 11589 2754 11627 2788
rect 11661 2754 11668 2788
rect 11476 2708 11668 2754
rect 11476 2674 11483 2708
rect 11517 2674 11555 2708
rect 11589 2674 11627 2708
rect 11661 2674 11668 2708
rect 11476 2657 11668 2674
rect 11476 2605 11482 2657
rect 11534 2605 11546 2657
rect 11598 2605 11610 2657
rect 11662 2605 11668 2657
rect 11476 2594 11483 2605
rect 11517 2594 11555 2605
rect 11589 2594 11627 2605
rect 11661 2594 11668 2605
rect 11476 2592 11668 2594
rect 11476 2540 11482 2592
rect 11534 2540 11546 2592
rect 11598 2540 11610 2592
rect 11662 2540 11668 2592
rect 11476 2527 11555 2540
rect 11589 2527 11668 2540
rect 11476 2475 11482 2527
rect 11534 2518 11546 2527
rect 11598 2518 11610 2527
rect 11662 2475 11668 2527
rect 11476 2462 11483 2475
rect 11661 2462 11668 2475
rect 11476 2410 11482 2462
rect 11662 2410 11668 2462
rect 11476 2397 11483 2410
rect 11661 2397 11668 2410
rect 11476 2345 11482 2397
rect 11662 2345 11668 2397
rect 11476 2332 11483 2345
rect 11661 2332 11668 2345
rect 11476 2280 11482 2332
rect 11662 2280 11668 2332
rect 11476 2267 11483 2280
rect 11661 2267 11668 2280
rect 11476 2215 11482 2267
rect 11662 2215 11668 2267
rect 11476 2202 11483 2215
rect 11661 2202 11668 2215
rect 11476 2150 11482 2202
rect 11662 2150 11668 2202
rect 11476 2137 11483 2150
rect 11661 2137 11668 2150
rect 11476 2085 11482 2137
rect 11662 2085 11668 2137
rect 11476 2072 11483 2085
rect 11661 2072 11668 2085
rect 11476 2020 11482 2072
rect 11662 2020 11668 2072
rect 11476 2007 11483 2020
rect 11661 2007 11668 2020
rect 11476 1955 11482 2007
rect 11662 1955 11668 2007
rect 11476 1942 11483 1955
rect 11661 1942 11668 1955
rect 11476 1890 11482 1942
rect 11662 1890 11668 1942
rect 11476 1877 11483 1890
rect 11661 1877 11668 1890
rect 11476 1825 11482 1877
rect 11662 1825 11668 1877
rect 11476 1812 11483 1825
rect 11661 1812 11668 1825
rect 11476 1568 11482 1812
rect 11662 1568 11668 1812
rect 11476 1562 11668 1568
rect 11972 4119 12164 4125
rect 11972 4067 11978 4119
rect 12030 4067 12042 4119
rect 12094 4067 12106 4119
rect 12158 4067 12164 4119
rect 11972 4064 11979 4067
rect 12013 4064 12051 4067
rect 12085 4064 12123 4067
rect 12157 4064 12164 4067
rect 11972 4054 12164 4064
rect 11972 4002 11978 4054
rect 12030 4002 12042 4054
rect 12094 4002 12106 4054
rect 12158 4002 12164 4054
rect 11972 3991 11979 4002
rect 12013 3991 12051 4002
rect 12085 3991 12123 4002
rect 12157 3991 12164 4002
rect 11972 3989 12164 3991
rect 11972 3937 11978 3989
rect 12030 3937 12042 3989
rect 12094 3937 12106 3989
rect 12158 3937 12164 3989
rect 11972 3924 11979 3937
rect 12013 3924 12051 3937
rect 12085 3924 12123 3937
rect 12157 3924 12164 3937
rect 11972 3872 11978 3924
rect 12030 3872 12042 3924
rect 12094 3872 12106 3924
rect 12158 3872 12164 3924
rect 11972 3859 11979 3872
rect 12013 3859 12051 3872
rect 12085 3859 12123 3872
rect 12157 3859 12164 3872
rect 11972 3807 11978 3859
rect 12030 3807 12042 3859
rect 12094 3807 12106 3859
rect 12158 3807 12164 3859
rect 11972 3806 12164 3807
rect 11972 3794 11979 3806
rect 12013 3794 12051 3806
rect 12085 3794 12123 3806
rect 12157 3794 12164 3806
rect 11972 3742 11978 3794
rect 12030 3742 12042 3794
rect 12094 3742 12106 3794
rect 12158 3742 12164 3794
rect 11972 3733 12164 3742
rect 11972 3729 11979 3733
rect 12013 3729 12051 3733
rect 12085 3729 12123 3733
rect 12157 3729 12164 3733
rect 11972 3677 11978 3729
rect 12030 3677 12042 3729
rect 12094 3677 12106 3729
rect 12158 3677 12164 3729
rect 11972 3664 12164 3677
rect 11972 2972 11978 3664
rect 12158 2972 12164 3664
rect 11972 2969 11979 2972
rect 12013 2969 12051 2972
rect 12085 2969 12123 2972
rect 12157 2969 12164 2972
rect 11972 2930 12164 2969
rect 11972 2896 11979 2930
rect 12013 2896 12051 2930
rect 12085 2896 12123 2930
rect 12157 2896 12164 2930
rect 11972 2857 12164 2896
rect 11972 2823 11979 2857
rect 12013 2823 12051 2857
rect 12085 2823 12123 2857
rect 12157 2823 12164 2857
rect 11972 2784 12164 2823
rect 11972 2750 11979 2784
rect 12013 2750 12051 2784
rect 12085 2750 12123 2784
rect 12157 2750 12164 2784
rect 11972 2711 12164 2750
rect 11972 2677 11979 2711
rect 12013 2677 12051 2711
rect 12085 2677 12123 2711
rect 12157 2677 12164 2711
rect 11972 2638 12164 2677
rect 11972 2604 11979 2638
rect 12013 2604 12051 2638
rect 12085 2604 12123 2638
rect 12157 2604 12164 2638
rect 11972 2565 12164 2604
rect 11972 2531 11979 2565
rect 12013 2531 12051 2565
rect 12085 2531 12123 2565
rect 12157 2531 12164 2565
rect 11972 2492 12164 2531
rect 11972 2458 11979 2492
rect 12013 2458 12051 2492
rect 12085 2458 12123 2492
rect 12157 2458 12164 2492
rect 11972 2419 12164 2458
rect 11972 2385 11979 2419
rect 12013 2385 12051 2419
rect 12085 2385 12123 2419
rect 12157 2385 12164 2419
rect 11972 2346 12164 2385
rect 11972 2312 11979 2346
rect 12013 2312 12051 2346
rect 12085 2312 12123 2346
rect 12157 2312 12164 2346
rect 11972 2273 12164 2312
rect 11972 2239 11979 2273
rect 12013 2239 12051 2273
rect 12085 2239 12123 2273
rect 12157 2239 12164 2273
rect 11972 2200 12164 2239
rect 11972 2166 11979 2200
rect 12013 2166 12051 2200
rect 12085 2166 12123 2200
rect 12157 2166 12164 2200
rect 11972 2126 12164 2166
rect 11972 2092 11979 2126
rect 12013 2092 12051 2126
rect 12085 2092 12123 2126
rect 12157 2092 12164 2126
rect 11972 2052 12164 2092
rect 11972 2018 11979 2052
rect 12013 2018 12051 2052
rect 12085 2018 12123 2052
rect 12157 2018 12164 2052
rect 11972 1978 12164 2018
rect 11972 1944 11979 1978
rect 12013 1944 12051 1978
rect 12085 1944 12123 1978
rect 12157 1944 12164 1978
rect 11972 1904 12164 1944
rect 11972 1870 11979 1904
rect 12013 1870 12051 1904
rect 12085 1870 12123 1904
rect 12157 1870 12164 1904
rect 11972 1830 12164 1870
rect 11972 1796 11979 1830
rect 12013 1796 12051 1830
rect 12085 1796 12123 1830
rect 12157 1796 12164 1830
rect 11972 1756 12164 1796
rect 11972 1722 11979 1756
rect 12013 1722 12051 1756
rect 12085 1722 12123 1756
rect 12157 1722 12164 1756
rect 11972 1682 12164 1722
rect 11972 1648 11979 1682
rect 12013 1648 12051 1682
rect 12085 1648 12123 1682
rect 12157 1648 12164 1682
rect 11972 1608 12164 1648
rect 11972 1574 11979 1608
rect 12013 1574 12051 1608
rect 12085 1574 12123 1608
rect 12157 1574 12164 1608
rect 11972 1562 12164 1574
rect 12468 4118 12660 4130
rect 12468 4092 12547 4118
rect 12581 4092 12660 4118
rect 12468 3194 12475 4092
rect 12653 3194 12660 4092
rect 12468 3182 12660 3194
rect 12468 3148 12547 3182
rect 12581 3148 12660 3182
rect 12468 3108 12660 3148
rect 12468 3074 12475 3108
rect 12509 3074 12547 3108
rect 12581 3074 12619 3108
rect 12653 3074 12660 3108
rect 12468 3028 12660 3074
rect 12468 2994 12475 3028
rect 12509 2994 12547 3028
rect 12581 2994 12619 3028
rect 12653 2994 12660 3028
rect 12468 2948 12660 2994
rect 12468 2914 12475 2948
rect 12509 2914 12547 2948
rect 12581 2914 12619 2948
rect 12653 2914 12660 2948
rect 12468 2868 12660 2914
rect 12468 2834 12475 2868
rect 12509 2834 12547 2868
rect 12581 2834 12619 2868
rect 12653 2834 12660 2868
rect 12468 2788 12660 2834
rect 12468 2754 12475 2788
rect 12509 2754 12547 2788
rect 12581 2754 12619 2788
rect 12653 2754 12660 2788
rect 12468 2708 12660 2754
rect 12468 2674 12475 2708
rect 12509 2674 12547 2708
rect 12581 2674 12619 2708
rect 12653 2674 12660 2708
rect 12468 2657 12660 2674
rect 12468 2605 12474 2657
rect 12526 2605 12538 2657
rect 12590 2605 12602 2657
rect 12654 2605 12660 2657
rect 12468 2594 12475 2605
rect 12509 2594 12547 2605
rect 12581 2594 12619 2605
rect 12653 2594 12660 2605
rect 12468 2592 12660 2594
rect 12468 2540 12474 2592
rect 12526 2540 12538 2592
rect 12590 2540 12602 2592
rect 12654 2540 12660 2592
rect 12468 2527 12547 2540
rect 12581 2527 12660 2540
rect 12468 2475 12474 2527
rect 12526 2518 12538 2527
rect 12590 2518 12602 2527
rect 12654 2475 12660 2527
rect 12468 2462 12475 2475
rect 12653 2462 12660 2475
rect 12468 2410 12474 2462
rect 12654 2410 12660 2462
rect 12468 2397 12475 2410
rect 12653 2397 12660 2410
rect 12468 2345 12474 2397
rect 12654 2345 12660 2397
rect 12468 2332 12475 2345
rect 12653 2332 12660 2345
rect 12468 2280 12474 2332
rect 12654 2280 12660 2332
rect 12468 2267 12475 2280
rect 12653 2267 12660 2280
rect 12468 2215 12474 2267
rect 12654 2215 12660 2267
rect 12468 2202 12475 2215
rect 12653 2202 12660 2215
rect 12468 2150 12474 2202
rect 12654 2150 12660 2202
rect 12468 2137 12475 2150
rect 12653 2137 12660 2150
rect 12468 2085 12474 2137
rect 12654 2085 12660 2137
rect 12468 2072 12475 2085
rect 12653 2072 12660 2085
rect 12468 2020 12474 2072
rect 12654 2020 12660 2072
rect 12468 2007 12475 2020
rect 12653 2007 12660 2020
rect 12468 1955 12474 2007
rect 12654 1955 12660 2007
rect 12468 1942 12475 1955
rect 12653 1942 12660 1955
rect 12468 1890 12474 1942
rect 12654 1890 12660 1942
rect 12468 1877 12475 1890
rect 12653 1877 12660 1890
rect 12468 1825 12474 1877
rect 12654 1825 12660 1877
rect 12468 1812 12475 1825
rect 12653 1812 12660 1825
rect 12468 1568 12474 1812
rect 12654 1568 12660 1812
rect 12468 1562 12660 1568
rect 12964 4119 13156 4125
rect 12964 4067 12970 4119
rect 13022 4067 13034 4119
rect 13086 4067 13098 4119
rect 13150 4067 13156 4119
rect 12964 4064 12971 4067
rect 13005 4064 13043 4067
rect 13077 4064 13115 4067
rect 13149 4064 13156 4067
rect 12964 4054 13156 4064
rect 12964 4002 12970 4054
rect 13022 4002 13034 4054
rect 13086 4002 13098 4054
rect 13150 4002 13156 4054
rect 12964 3991 12971 4002
rect 13005 3991 13043 4002
rect 13077 3991 13115 4002
rect 13149 3991 13156 4002
rect 12964 3989 13156 3991
rect 12964 3937 12970 3989
rect 13022 3937 13034 3989
rect 13086 3937 13098 3989
rect 13150 3937 13156 3989
rect 12964 3924 12971 3937
rect 13005 3924 13043 3937
rect 13077 3924 13115 3937
rect 13149 3924 13156 3937
rect 12964 3872 12970 3924
rect 13022 3872 13034 3924
rect 13086 3872 13098 3924
rect 13150 3872 13156 3924
rect 12964 3859 12971 3872
rect 13005 3859 13043 3872
rect 13077 3859 13115 3872
rect 13149 3859 13156 3872
rect 12964 3807 12970 3859
rect 13022 3807 13034 3859
rect 13086 3807 13098 3859
rect 13150 3807 13156 3859
rect 12964 3806 13156 3807
rect 12964 3794 12971 3806
rect 13005 3794 13043 3806
rect 13077 3794 13115 3806
rect 13149 3794 13156 3806
rect 12964 3742 12970 3794
rect 13022 3742 13034 3794
rect 13086 3742 13098 3794
rect 13150 3742 13156 3794
rect 12964 3733 13156 3742
rect 12964 3729 12971 3733
rect 13005 3729 13043 3733
rect 13077 3729 13115 3733
rect 13149 3729 13156 3733
rect 12964 3677 12970 3729
rect 13022 3677 13034 3729
rect 13086 3677 13098 3729
rect 13150 3677 13156 3729
rect 12964 3664 13156 3677
rect 12964 2972 12970 3664
rect 13150 2972 13156 3664
rect 12964 2969 12971 2972
rect 13005 2969 13043 2972
rect 13077 2969 13115 2972
rect 13149 2969 13156 2972
rect 12964 2930 13156 2969
rect 12964 2896 12971 2930
rect 13005 2896 13043 2930
rect 13077 2896 13115 2930
rect 13149 2896 13156 2930
rect 12964 2857 13156 2896
rect 12964 2823 12971 2857
rect 13005 2823 13043 2857
rect 13077 2823 13115 2857
rect 13149 2823 13156 2857
rect 12964 2784 13156 2823
rect 12964 2750 12971 2784
rect 13005 2750 13043 2784
rect 13077 2750 13115 2784
rect 13149 2750 13156 2784
rect 12964 2711 13156 2750
rect 12964 2677 12971 2711
rect 13005 2677 13043 2711
rect 13077 2677 13115 2711
rect 13149 2677 13156 2711
rect 12964 2638 13156 2677
rect 12964 2604 12971 2638
rect 13005 2604 13043 2638
rect 13077 2604 13115 2638
rect 13149 2604 13156 2638
rect 12964 2565 13156 2604
rect 12964 2531 12971 2565
rect 13005 2531 13043 2565
rect 13077 2531 13115 2565
rect 13149 2531 13156 2565
rect 12964 2492 13156 2531
rect 12964 2458 12971 2492
rect 13005 2458 13043 2492
rect 13077 2458 13115 2492
rect 13149 2458 13156 2492
rect 12964 2419 13156 2458
rect 12964 2385 12971 2419
rect 13005 2385 13043 2419
rect 13077 2385 13115 2419
rect 13149 2385 13156 2419
rect 12964 2346 13156 2385
rect 12964 2312 12971 2346
rect 13005 2312 13043 2346
rect 13077 2312 13115 2346
rect 13149 2312 13156 2346
rect 12964 2273 13156 2312
rect 12964 2239 12971 2273
rect 13005 2239 13043 2273
rect 13077 2239 13115 2273
rect 13149 2239 13156 2273
rect 12964 2200 13156 2239
rect 12964 2166 12971 2200
rect 13005 2166 13043 2200
rect 13077 2166 13115 2200
rect 13149 2166 13156 2200
rect 12964 2126 13156 2166
rect 12964 2092 12971 2126
rect 13005 2092 13043 2126
rect 13077 2092 13115 2126
rect 13149 2092 13156 2126
rect 12964 2052 13156 2092
rect 12964 2018 12971 2052
rect 13005 2018 13043 2052
rect 13077 2018 13115 2052
rect 13149 2018 13156 2052
rect 12964 1978 13156 2018
rect 12964 1944 12971 1978
rect 13005 1944 13043 1978
rect 13077 1944 13115 1978
rect 13149 1944 13156 1978
rect 12964 1904 13156 1944
rect 12964 1870 12971 1904
rect 13005 1870 13043 1904
rect 13077 1870 13115 1904
rect 13149 1870 13156 1904
rect 12964 1830 13156 1870
rect 12964 1796 12971 1830
rect 13005 1796 13043 1830
rect 13077 1796 13115 1830
rect 13149 1796 13156 1830
rect 12964 1756 13156 1796
rect 12964 1722 12971 1756
rect 13005 1722 13043 1756
rect 13077 1722 13115 1756
rect 13149 1722 13156 1756
rect 12964 1682 13156 1722
rect 12964 1648 12971 1682
rect 13005 1648 13043 1682
rect 13077 1648 13115 1682
rect 13149 1648 13156 1682
rect 12964 1608 13156 1648
rect 12964 1574 12971 1608
rect 13005 1574 13043 1608
rect 13077 1574 13115 1608
rect 13149 1574 13156 1608
rect 12964 1562 13156 1574
rect 13460 4118 13652 4130
rect 13460 4092 13539 4118
rect 13573 4092 13652 4118
rect 13460 3194 13467 4092
rect 13645 3194 13652 4092
rect 13460 3182 13652 3194
rect 13460 3148 13539 3182
rect 13573 3148 13652 3182
rect 13460 3108 13652 3148
rect 13460 3074 13467 3108
rect 13501 3074 13539 3108
rect 13573 3074 13611 3108
rect 13645 3074 13652 3108
rect 13460 3028 13652 3074
rect 13460 2994 13467 3028
rect 13501 2994 13539 3028
rect 13573 2994 13611 3028
rect 13645 2994 13652 3028
rect 13460 2948 13652 2994
rect 13460 2914 13467 2948
rect 13501 2914 13539 2948
rect 13573 2914 13611 2948
rect 13645 2914 13652 2948
rect 13460 2868 13652 2914
rect 13460 2834 13467 2868
rect 13501 2834 13539 2868
rect 13573 2834 13611 2868
rect 13645 2834 13652 2868
rect 13460 2788 13652 2834
rect 13460 2754 13467 2788
rect 13501 2754 13539 2788
rect 13573 2754 13611 2788
rect 13645 2754 13652 2788
rect 13460 2708 13652 2754
rect 13460 2674 13467 2708
rect 13501 2674 13539 2708
rect 13573 2674 13611 2708
rect 13645 2674 13652 2708
rect 13460 2657 13652 2674
rect 13460 2605 13466 2657
rect 13518 2605 13530 2657
rect 13582 2605 13594 2657
rect 13646 2605 13652 2657
rect 13460 2594 13467 2605
rect 13501 2594 13539 2605
rect 13573 2594 13611 2605
rect 13645 2594 13652 2605
rect 13460 2592 13652 2594
rect 13460 2540 13466 2592
rect 13518 2540 13530 2592
rect 13582 2540 13594 2592
rect 13646 2540 13652 2592
rect 13460 2527 13539 2540
rect 13573 2527 13652 2540
rect 13460 2475 13466 2527
rect 13518 2518 13530 2527
rect 13582 2518 13594 2527
rect 13646 2475 13652 2527
rect 13460 2462 13467 2475
rect 13645 2462 13652 2475
rect 13460 2410 13466 2462
rect 13646 2410 13652 2462
rect 13460 2397 13467 2410
rect 13645 2397 13652 2410
rect 13460 2345 13466 2397
rect 13646 2345 13652 2397
rect 13460 2332 13467 2345
rect 13645 2332 13652 2345
rect 13460 2280 13466 2332
rect 13646 2280 13652 2332
rect 13460 2267 13467 2280
rect 13645 2267 13652 2280
rect 13460 2215 13466 2267
rect 13646 2215 13652 2267
rect 13460 2202 13467 2215
rect 13645 2202 13652 2215
rect 13460 2150 13466 2202
rect 13646 2150 13652 2202
rect 13460 2137 13467 2150
rect 13645 2137 13652 2150
rect 13460 2085 13466 2137
rect 13646 2085 13652 2137
rect 13460 2072 13467 2085
rect 13645 2072 13652 2085
rect 13460 2020 13466 2072
rect 13646 2020 13652 2072
rect 13460 2007 13467 2020
rect 13645 2007 13652 2020
rect 13460 1955 13466 2007
rect 13646 1955 13652 2007
rect 13460 1942 13467 1955
rect 13645 1942 13652 1955
rect 13460 1890 13466 1942
rect 13646 1890 13652 1942
rect 13460 1877 13467 1890
rect 13645 1877 13652 1890
rect 13460 1825 13466 1877
rect 13646 1825 13652 1877
rect 13460 1812 13467 1825
rect 13645 1812 13652 1825
rect 13460 1568 13466 1812
rect 13646 1568 13652 1812
rect 13460 1562 13652 1568
rect 13990 4119 14135 4130
rect 14042 4067 14062 4119
rect 14114 4067 14135 4119
rect 13990 4064 13999 4067
rect 14033 4064 14135 4067
rect 13990 4055 14135 4064
rect 14042 4003 14062 4055
rect 14114 4003 14135 4055
rect 13990 3991 13999 4003
rect 14033 3991 14135 4003
rect 14042 3939 14062 3991
rect 14114 3939 14135 3991
rect 13990 3927 13999 3939
rect 14033 3927 14135 3939
rect 14042 3875 14062 3927
rect 14114 3875 14135 3927
rect 13990 3863 13999 3875
rect 14033 3863 14135 3875
rect 14042 3811 14062 3863
rect 14114 3811 14135 3863
rect 13990 3806 14135 3811
rect 13990 3799 13999 3806
rect 14033 3799 14135 3806
rect 14042 3747 14062 3799
rect 14114 3747 14135 3799
rect 13990 3735 14135 3747
rect 14042 3683 14062 3735
rect 14114 3683 14135 3735
rect 13990 3671 14135 3683
rect 14042 3619 14062 3671
rect 14114 3619 14135 3671
rect 13990 3607 14135 3619
rect 14042 3555 14062 3607
rect 14114 3555 14135 3607
rect 13990 3553 13999 3555
rect 14033 3553 14135 3555
rect 13990 3543 14135 3553
rect 14042 3491 14062 3543
rect 14114 3491 14135 3543
rect 13990 3480 13999 3491
rect 14033 3480 14135 3491
rect 13990 3479 14135 3480
rect 14042 3427 14062 3479
rect 14114 3427 14135 3479
rect 13990 3414 13999 3427
rect 14033 3414 14135 3427
rect 14042 3362 14062 3414
rect 14114 3362 14135 3414
rect 13990 3349 13999 3362
rect 14033 3349 14135 3362
rect 14042 3297 14062 3349
rect 14114 3297 14135 3349
rect 13990 3295 14135 3297
rect 13990 3284 13999 3295
rect 14033 3284 14135 3295
rect 14042 3232 14062 3284
rect 14114 3232 14135 3284
rect 13990 3222 14135 3232
rect 13990 3219 13999 3222
rect 14033 3219 14135 3222
rect 14042 3167 14062 3219
rect 14114 3167 14135 3219
rect 13990 3154 14135 3167
rect 14042 3102 14062 3154
rect 14114 3102 14135 3154
rect 13990 3089 14135 3102
rect 14042 3037 14062 3089
rect 14114 3037 14135 3089
rect 13990 3024 14135 3037
rect 14042 2972 14062 3024
rect 14114 2972 14135 3024
rect 13990 2969 13999 2972
rect 14033 2969 14135 2972
rect 13990 2930 14135 2969
rect 13990 2896 13999 2930
rect 14033 2896 14135 2930
rect 13990 2857 14135 2896
rect 13990 2823 13999 2857
rect 14033 2823 14135 2857
rect 13990 2784 14135 2823
rect 13990 2750 13999 2784
rect 14033 2750 14135 2784
rect 13990 2711 14135 2750
rect 13990 2677 13999 2711
rect 14033 2677 14135 2711
rect 13990 2638 14135 2677
rect 13990 2604 13999 2638
rect 14033 2604 14135 2638
rect 13990 2565 14135 2604
rect 13990 2531 13999 2565
rect 14033 2531 14135 2565
rect 13990 2492 14135 2531
rect 13990 2458 13999 2492
rect 14033 2458 14135 2492
rect 13990 2419 14135 2458
rect 13990 2385 13999 2419
rect 14033 2385 14135 2419
rect 13990 2346 14135 2385
rect 13990 2312 13999 2346
rect 14033 2312 14135 2346
rect 13990 2273 14135 2312
rect 13990 2239 13999 2273
rect 14033 2239 14135 2273
rect 13990 2200 14135 2239
rect 13990 2166 13999 2200
rect 14033 2166 14135 2200
rect 13990 2126 14135 2166
rect 13990 2092 13999 2126
rect 14033 2092 14135 2126
rect 13990 2052 14135 2092
rect 13990 2018 13999 2052
rect 14033 2018 14135 2052
rect 13990 1978 14135 2018
rect 13990 1944 13999 1978
rect 14033 1944 14135 1978
rect 13990 1904 14135 1944
rect 13990 1870 13999 1904
rect 14033 1870 14135 1904
rect 13990 1830 14135 1870
rect 13990 1796 13999 1830
rect 14033 1796 14135 1830
rect 13990 1756 14135 1796
rect 13990 1722 13999 1756
rect 14033 1722 14135 1756
rect 13990 1682 14135 1722
rect 13990 1648 13999 1682
rect 14033 1648 14135 1682
rect 13990 1608 14135 1648
rect 13990 1574 13999 1608
rect 14033 1574 14135 1608
rect 13990 1536 14135 1574
rect 14350 4106 14356 4140
rect 14390 4106 14428 4140
rect 14350 4067 14428 4106
rect 14350 4033 14356 4067
rect 14390 4033 14428 4067
rect 14350 3994 14428 4033
rect 14350 3960 14356 3994
rect 14390 3960 14428 3994
rect 14606 3960 14618 4426
rect 14350 3952 14618 3960
rect 14350 3921 14428 3952
rect 14350 3887 14356 3921
rect 14390 3918 14428 3921
rect 14462 3921 14618 3952
rect 14462 3918 14500 3921
rect 14390 3887 14500 3918
rect 14534 3887 14572 3921
rect 14606 3887 14618 3921
rect 14350 3880 14618 3887
rect 14350 3848 14428 3880
rect 14350 3814 14356 3848
rect 14390 3846 14428 3848
rect 14462 3848 14618 3880
rect 14462 3846 14500 3848
rect 14390 3814 14500 3846
rect 14534 3814 14572 3848
rect 14606 3814 14618 3848
rect 14350 3808 14618 3814
rect 14350 3775 14428 3808
rect 14350 3741 14356 3775
rect 14390 3774 14428 3775
rect 14462 3775 14618 3808
rect 14462 3774 14500 3775
rect 14390 3741 14500 3774
rect 14534 3741 14572 3775
rect 14606 3741 14618 3775
rect 14350 3736 14618 3741
rect 14350 3702 14428 3736
rect 14462 3702 14618 3736
rect 14350 3668 14356 3702
rect 14390 3668 14500 3702
rect 14534 3668 14572 3702
rect 14606 3668 14618 3702
rect 14350 3664 14618 3668
rect 14350 3630 14428 3664
rect 14462 3630 14618 3664
rect 14350 3629 14618 3630
rect 14350 3595 14356 3629
rect 14390 3595 14500 3629
rect 14534 3595 14572 3629
rect 14606 3595 14618 3629
rect 14350 3592 14618 3595
rect 14350 3558 14428 3592
rect 14462 3558 14618 3592
rect 14350 3556 14618 3558
rect 14350 3522 14356 3556
rect 14390 3522 14500 3556
rect 14534 3522 14572 3556
rect 14606 3522 14618 3556
rect 14350 3520 14618 3522
rect 14350 3486 14428 3520
rect 14462 3486 14618 3520
rect 14350 3483 14618 3486
rect 14350 3449 14356 3483
rect 14390 3449 14500 3483
rect 14534 3449 14572 3483
rect 14606 3449 14618 3483
rect 14350 3448 14618 3449
rect 14350 3414 14428 3448
rect 14462 3414 14618 3448
rect 14350 3410 14618 3414
rect 14350 3376 14356 3410
rect 14390 3376 14500 3410
rect 14534 3376 14572 3410
rect 14606 3376 14618 3410
rect 14350 3342 14428 3376
rect 14462 3342 14618 3376
rect 14350 3337 14618 3342
rect 14350 3303 14356 3337
rect 14390 3304 14500 3337
rect 14390 3303 14428 3304
rect 14350 3270 14428 3303
rect 14462 3303 14500 3304
rect 14534 3303 14572 3337
rect 14606 3303 14618 3337
rect 14462 3270 14618 3303
rect 14350 3264 14618 3270
rect 14350 3230 14356 3264
rect 14390 3232 14500 3264
rect 14390 3230 14428 3232
rect 14350 3198 14428 3230
rect 14462 3230 14500 3232
rect 14534 3230 14572 3264
rect 14606 3230 14618 3264
rect 14462 3198 14618 3230
rect 14350 3191 14618 3198
rect 14350 3157 14356 3191
rect 14390 3160 14500 3191
rect 14390 3157 14428 3160
rect 14350 3126 14428 3157
rect 14462 3157 14500 3160
rect 14534 3157 14572 3191
rect 14606 3157 14618 3191
rect 14462 3126 14618 3157
rect 14350 3118 14618 3126
rect 14350 3084 14356 3118
rect 14390 3088 14500 3118
rect 14390 3084 14428 3088
rect 14350 3054 14428 3084
rect 14462 3084 14500 3088
rect 14534 3084 14572 3118
rect 14606 3084 14618 3118
rect 14462 3054 14618 3084
rect 14350 3045 14618 3054
rect 14350 3011 14356 3045
rect 14390 3016 14500 3045
rect 14390 3011 14428 3016
rect 14350 2982 14428 3011
rect 14462 3011 14500 3016
rect 14534 3011 14572 3045
rect 14606 3011 14618 3045
rect 14462 2982 14618 3011
rect 14350 2972 14618 2982
rect 14350 2938 14356 2972
rect 14390 2944 14500 2972
rect 14390 2938 14428 2944
rect 14350 2910 14428 2938
rect 14462 2938 14500 2944
rect 14534 2938 14572 2972
rect 14606 2938 14618 2972
rect 14462 2910 14618 2938
rect 14350 2899 14618 2910
rect 14350 2865 14356 2899
rect 14390 2872 14500 2899
rect 14390 2865 14428 2872
rect 14350 2838 14428 2865
rect 14462 2865 14500 2872
rect 14534 2865 14572 2899
rect 14606 2865 14618 2899
rect 14462 2838 14618 2865
rect 14350 2826 14618 2838
rect 14350 2792 14356 2826
rect 14390 2800 14500 2826
rect 14390 2792 14428 2800
rect 14350 2766 14428 2792
rect 14462 2792 14500 2800
rect 14534 2792 14572 2826
rect 14606 2792 14618 2826
rect 14462 2766 14618 2792
rect 14350 2753 14618 2766
rect 14350 2719 14356 2753
rect 14390 2728 14500 2753
rect 14390 2719 14428 2728
rect 14350 2694 14428 2719
rect 14462 2719 14500 2728
rect 14534 2719 14572 2753
rect 14606 2719 14618 2753
rect 14462 2694 14618 2719
rect 14350 2680 14618 2694
rect 14350 2657 14356 2680
rect 14390 2657 14500 2680
rect 14534 2657 14572 2680
rect 14606 2657 14618 2680
rect 14402 2605 14422 2657
rect 14474 2605 14494 2657
rect 14546 2605 14566 2657
rect 14350 2592 14356 2605
rect 14390 2592 14500 2605
rect 14534 2592 14572 2605
rect 14606 2592 14618 2605
rect 14402 2540 14422 2592
rect 14474 2540 14494 2592
rect 14546 2540 14566 2592
rect 14350 2534 14618 2540
rect 14350 2527 14356 2534
rect 14390 2527 14500 2534
rect 14534 2527 14572 2534
rect 14606 2527 14618 2534
rect 14402 2475 14422 2527
rect 14474 2475 14494 2527
rect 14546 2475 14566 2527
rect 14350 2462 14618 2475
rect 14402 2410 14422 2462
rect 14474 2410 14494 2462
rect 14546 2410 14566 2462
rect 14350 2406 14428 2410
rect 14462 2406 14618 2410
rect 14350 2397 14618 2406
rect 14402 2345 14422 2397
rect 14474 2345 14494 2397
rect 14546 2345 14566 2397
rect 14350 2334 14428 2345
rect 14462 2334 14618 2345
rect 14350 2332 14618 2334
rect 14402 2280 14422 2332
rect 14474 2280 14494 2332
rect 14546 2280 14566 2332
rect 14350 2267 14428 2280
rect 14462 2267 14618 2280
rect 14402 2215 14422 2267
rect 14474 2215 14494 2267
rect 14546 2215 14566 2267
rect 14350 2208 14356 2215
rect 14390 2208 14428 2215
rect 14350 2202 14428 2208
rect 14462 2208 14500 2215
rect 14534 2208 14572 2215
rect 14606 2208 14618 2215
rect 14462 2202 14618 2208
rect 14402 2150 14422 2202
rect 14474 2150 14494 2202
rect 14546 2150 14566 2202
rect 14350 2137 14356 2150
rect 14390 2137 14428 2150
rect 14462 2137 14500 2150
rect 14534 2137 14572 2150
rect 14606 2137 14618 2150
rect 14402 2085 14422 2137
rect 14474 2085 14494 2137
rect 14546 2085 14566 2137
rect 14350 2072 14356 2085
rect 14390 2080 14500 2085
rect 14390 2072 14428 2080
rect 14462 2072 14500 2080
rect 14534 2072 14572 2085
rect 14606 2072 14618 2085
rect 14402 2020 14422 2072
rect 14474 2020 14494 2072
rect 14546 2020 14566 2072
rect 14350 2007 14356 2020
rect 14390 2008 14500 2020
rect 14390 2007 14428 2008
rect 14462 2007 14500 2008
rect 14534 2007 14572 2020
rect 14606 2007 14618 2020
rect 14402 1955 14422 2007
rect 14474 1955 14494 2007
rect 14546 1955 14566 2007
rect 14350 1950 14618 1955
rect 14350 1942 14356 1950
rect 14390 1942 14500 1950
rect 14534 1942 14572 1950
rect 14606 1942 14618 1950
rect 14402 1890 14422 1942
rect 14474 1890 14494 1942
rect 14546 1890 14566 1942
rect 14350 1877 14618 1890
rect 14402 1825 14422 1877
rect 14474 1825 14494 1877
rect 14546 1825 14566 1877
rect 14350 1812 14618 1825
rect 14402 1760 14422 1812
rect 14474 1760 14494 1812
rect 14546 1760 14566 1812
rect 14350 1758 14428 1760
rect 14462 1758 14618 1760
rect 14350 1748 14618 1758
rect 14402 1696 14422 1748
rect 14474 1696 14494 1748
rect 14546 1696 14566 1748
rect 14350 1686 14428 1696
rect 14462 1686 14618 1696
rect 14350 1684 14618 1686
rect 14402 1632 14422 1684
rect 14474 1632 14494 1684
rect 14546 1632 14566 1684
rect 14350 1623 14356 1632
rect 14390 1623 14428 1632
rect 14350 1620 14428 1623
rect 14462 1624 14500 1632
rect 14534 1624 14572 1632
rect 14606 1624 14618 1632
rect 14462 1620 14618 1624
rect 14402 1568 14422 1620
rect 14474 1568 14494 1620
rect 14546 1568 14566 1620
rect 14350 1549 14356 1568
rect 14390 1549 14428 1568
rect 14350 1542 14428 1549
rect 14462 1551 14500 1568
rect 14534 1551 14572 1568
rect 14606 1551 14618 1568
rect 14462 1542 14618 1551
rect 14350 1512 14618 1542
rect 14350 1509 14500 1512
rect 14350 1475 14356 1509
rect 14390 1504 14500 1509
rect 14390 1475 14428 1504
rect 14350 1470 14428 1475
rect 14462 1478 14500 1504
rect 14534 1478 14572 1512
rect 14606 1478 14618 1512
rect 14462 1470 14618 1478
rect 14350 1439 14618 1470
rect 14350 1435 14500 1439
rect 14350 1401 14356 1435
rect 14390 1432 14500 1435
rect 14390 1401 14428 1432
rect 14350 1398 14428 1401
rect 14462 1405 14500 1432
rect 14534 1405 14572 1439
rect 14606 1405 14618 1439
rect 14462 1398 14618 1405
rect 14350 1366 14618 1398
rect 14350 1361 14500 1366
rect 14350 1327 14356 1361
rect 14390 1360 14500 1361
rect 14390 1327 14428 1360
rect 14350 1326 14428 1327
rect 14462 1332 14500 1360
rect 14534 1332 14572 1366
rect 14606 1332 14618 1366
rect 14462 1326 14618 1332
rect 14350 1293 14618 1326
rect 14350 1288 14500 1293
rect 14350 1287 14428 1288
rect 912 1250 970 1262
rect 912 1216 924 1250
rect 958 1216 970 1250
rect 912 1178 970 1216
rect 912 1144 924 1178
rect 958 1144 970 1178
rect 912 1132 970 1144
rect 1306 1250 1436 1262
rect 1306 1144 1318 1250
rect 1424 1144 1436 1250
rect 1306 1132 1436 1144
rect 1868 1250 1998 1262
rect 1868 1144 1880 1250
rect 1986 1144 1998 1250
rect 1868 1132 1998 1144
rect 2298 1250 2428 1262
rect 2298 1144 2310 1250
rect 2416 1144 2428 1250
rect 2298 1132 2428 1144
rect 2860 1250 2990 1262
rect 2860 1144 2872 1250
rect 2978 1144 2990 1250
rect 2860 1132 2990 1144
rect 3290 1250 3420 1262
rect 3290 1144 3302 1250
rect 3408 1144 3420 1250
rect 3290 1132 3420 1144
rect 3852 1250 3982 1262
rect 3852 1144 3864 1250
rect 3970 1144 3982 1250
rect 3852 1132 3982 1144
rect 4282 1250 4412 1262
rect 4282 1144 4294 1250
rect 4400 1144 4412 1250
rect 4282 1132 4412 1144
rect 4844 1250 4974 1262
rect 4844 1144 4856 1250
rect 4962 1144 4974 1250
rect 4844 1132 4974 1144
rect 5274 1250 5404 1262
rect 5274 1144 5286 1250
rect 5392 1144 5404 1250
rect 5274 1132 5404 1144
rect 5836 1250 5966 1262
rect 5836 1144 5848 1250
rect 5954 1144 5966 1250
rect 5836 1132 5966 1144
rect 6266 1250 6396 1262
rect 6266 1144 6278 1250
rect 6384 1144 6396 1250
rect 6266 1132 6396 1144
rect 6828 1250 6958 1262
rect 6828 1144 6840 1250
rect 6946 1144 6958 1250
rect 6828 1132 6958 1144
rect 7258 1250 7388 1262
rect 7258 1144 7270 1250
rect 7376 1144 7388 1250
rect 7258 1132 7388 1144
rect 7820 1250 7950 1262
rect 7820 1144 7832 1250
rect 7938 1144 7950 1250
rect 7820 1132 7950 1144
rect 8250 1250 8380 1262
rect 8250 1144 8262 1250
rect 8368 1144 8380 1250
rect 8250 1132 8380 1144
rect 8812 1250 8942 1262
rect 8812 1144 8824 1250
rect 8930 1144 8942 1250
rect 8812 1132 8942 1144
rect 9242 1250 9372 1262
rect 9242 1144 9254 1250
rect 9360 1144 9372 1250
rect 9242 1132 9372 1144
rect 9804 1250 9934 1262
rect 9804 1144 9816 1250
rect 9922 1144 9934 1250
rect 9804 1132 9934 1144
rect 10234 1250 10364 1262
rect 10234 1144 10246 1250
rect 10352 1144 10364 1250
rect 10234 1132 10364 1144
rect 10796 1250 10926 1262
rect 10796 1144 10808 1250
rect 10914 1144 10926 1250
rect 10796 1132 10926 1144
rect 11226 1250 11356 1262
rect 11226 1144 11238 1250
rect 11344 1144 11356 1250
rect 11226 1132 11356 1144
rect 11788 1250 11918 1262
rect 11788 1144 11800 1250
rect 11906 1144 11918 1250
rect 11788 1132 11918 1144
rect 12218 1250 12348 1262
rect 12218 1144 12230 1250
rect 12336 1144 12348 1250
rect 12218 1132 12348 1144
rect 12780 1250 12910 1262
rect 12780 1144 12792 1250
rect 12898 1144 12910 1250
rect 12780 1132 12910 1144
rect 13210 1250 13340 1262
rect 13210 1144 13222 1250
rect 13328 1144 13340 1250
rect 13210 1132 13340 1144
rect 13772 1250 13902 1262
rect 13772 1144 13784 1250
rect 13890 1144 13902 1250
rect 13772 1132 13902 1144
rect 14130 1250 14260 1262
rect 14130 1144 14142 1250
rect 14248 1144 14260 1250
rect 14130 1132 14260 1144
rect 14350 1253 14356 1287
rect 14390 1254 14428 1287
rect 14462 1259 14500 1288
rect 14534 1259 14572 1293
rect 14606 1259 14618 1293
rect 14462 1254 14618 1259
rect 14390 1253 14618 1254
rect 14350 1220 14618 1253
rect 14350 1216 14500 1220
rect 14350 1213 14428 1216
rect 14350 1179 14356 1213
rect 14390 1182 14428 1213
rect 14462 1186 14500 1216
rect 14534 1186 14572 1220
rect 14606 1186 14618 1220
rect 14462 1182 14618 1186
rect 14390 1179 14618 1182
rect 14350 1147 14618 1179
rect 14350 1144 14500 1147
rect 14350 1139 14428 1144
rect 14350 1105 14356 1139
rect 14390 1110 14428 1139
rect 14462 1113 14500 1144
rect 14534 1113 14572 1147
rect 14606 1113 14618 1147
rect 14462 1110 14618 1113
rect 14390 1105 14618 1110
rect 14350 1074 14618 1105
rect 14350 1072 14500 1074
rect 14350 1065 14428 1072
rect 14350 1031 14356 1065
rect 14390 1038 14428 1065
rect 14462 1040 14500 1072
rect 14534 1040 14572 1074
rect 14606 1040 14618 1074
rect 14462 1038 14618 1040
rect 14390 1031 14618 1038
tri 14349 1024 14350 1025 se
rect 14350 1024 14618 1031
tri 786 1001 809 1024 sw
tri 14326 1001 14349 1024 se
rect 14349 1001 14618 1024
rect 780 1000 809 1001
tri 809 1000 810 1001 sw
tri 14325 1000 14326 1001 se
rect 14326 1000 14500 1001
rect 780 991 810 1000
tri 810 991 819 1000 sw
tri 14316 991 14325 1000 se
rect 14325 991 14428 1000
rect 780 957 819 991
tri 819 957 853 991 sw
tri 14282 957 14316 991 se
rect 14316 957 14356 991
rect 14390 966 14428 991
rect 14462 967 14500 1000
rect 14534 967 14572 1001
rect 14606 967 14618 1001
rect 14462 966 14618 967
rect 14390 957 14618 966
rect 780 928 853 957
tri 853 928 882 957 sw
tri 14253 928 14282 957 se
rect 14282 928 14618 957
rect 780 917 882 928
tri 882 917 893 928 sw
tri 14242 917 14253 928 se
rect 14253 917 14428 928
rect 517 883 746 894
rect 780 883 893 917
tri 893 883 927 917 sw
tri 14208 883 14242 917 se
rect 14242 883 14356 917
rect 14390 894 14428 917
rect 14462 894 14500 928
rect 14534 894 14572 928
rect 14606 894 14618 928
rect 14390 883 14618 894
rect 229 829 269 863
rect 303 845 329 863
tri 329 845 366 882 sw
rect 517 872 927 883
tri 927 872 938 883 sw
tri 14197 872 14208 883 se
rect 14208 872 14618 883
rect 517 845 938 872
tri 938 845 965 872 sw
tri 14196 871 14197 872 se
rect 14197 871 14618 872
tri 14184 859 14196 871 se
rect 14196 859 14618 871
rect 14807 4420 14832 4454
rect 14866 4420 14907 4454
rect 14807 4382 14907 4420
rect 14807 4348 14832 4382
rect 14866 4348 14907 4382
rect 14807 4310 14907 4348
rect 14807 4276 14832 4310
rect 14866 4276 14907 4310
rect 14807 4238 14907 4276
rect 14807 4204 14832 4238
rect 14866 4204 14907 4238
rect 14807 4166 14907 4204
rect 14807 4132 14832 4166
rect 14866 4132 14907 4166
rect 14807 4094 14907 4132
rect 14807 4060 14832 4094
rect 14866 4060 14907 4094
rect 14807 4022 14907 4060
rect 14807 3988 14832 4022
rect 14866 3988 14907 4022
rect 14807 3950 14907 3988
rect 14807 3916 14832 3950
rect 14866 3916 14907 3950
rect 14807 3878 14907 3916
rect 14807 3844 14832 3878
rect 14866 3844 14907 3878
rect 14807 3806 14907 3844
rect 14807 3772 14832 3806
rect 14866 3772 14907 3806
rect 14807 3734 14907 3772
rect 14807 3700 14832 3734
rect 14866 3700 14907 3734
rect 14807 3662 14907 3700
rect 14807 3628 14832 3662
rect 14866 3628 14907 3662
rect 14807 3590 14907 3628
rect 14807 3556 14832 3590
rect 14866 3556 14907 3590
rect 14807 3518 14907 3556
rect 14807 3484 14832 3518
rect 14866 3484 14907 3518
rect 14807 3446 14907 3484
rect 14807 3412 14832 3446
rect 14866 3412 14907 3446
rect 14807 3374 14907 3412
rect 14807 3340 14832 3374
rect 14866 3340 14907 3374
rect 14807 3302 14907 3340
rect 14807 3268 14832 3302
rect 14866 3268 14907 3302
rect 14807 3230 14907 3268
rect 14807 3196 14832 3230
rect 14866 3196 14907 3230
rect 14807 3158 14907 3196
rect 14807 3124 14832 3158
rect 14866 3124 14907 3158
rect 14807 3086 14907 3124
rect 14807 3052 14832 3086
rect 14866 3052 14907 3086
rect 14807 3014 14907 3052
rect 14807 2980 14832 3014
rect 14866 2980 14907 3014
rect 14807 2942 14907 2980
rect 14807 2908 14832 2942
rect 14866 2908 14907 2942
rect 14807 2870 14907 2908
rect 14807 2836 14832 2870
rect 14866 2836 14907 2870
rect 14807 2798 14907 2836
rect 14807 2764 14832 2798
rect 14866 2764 14907 2798
rect 14807 2726 14907 2764
rect 14807 2692 14832 2726
rect 14866 2692 14907 2726
rect 14807 2654 14907 2692
rect 14807 2620 14832 2654
rect 14866 2620 14907 2654
rect 14807 2582 14907 2620
rect 14807 2548 14832 2582
rect 14866 2548 14907 2582
rect 14807 2510 14907 2548
rect 14807 2476 14832 2510
rect 14866 2476 14907 2510
rect 14807 2438 14907 2476
rect 14807 2404 14832 2438
rect 14866 2404 14907 2438
rect 14807 2366 14907 2404
rect 14807 2332 14832 2366
rect 14866 2332 14907 2366
rect 14807 2294 14907 2332
rect 14807 2260 14832 2294
rect 14866 2260 14907 2294
rect 14807 2222 14907 2260
rect 14807 2188 14832 2222
rect 14866 2188 14907 2222
rect 14807 2150 14907 2188
rect 14807 2116 14832 2150
rect 14866 2116 14907 2150
rect 14807 2078 14907 2116
rect 14807 2044 14832 2078
rect 14866 2044 14907 2078
rect 14807 2006 14907 2044
rect 14807 1972 14832 2006
rect 14866 1972 14907 2006
rect 14807 1934 14907 1972
rect 14807 1900 14832 1934
rect 14866 1900 14907 1934
rect 14807 1862 14907 1900
rect 14807 1828 14832 1862
rect 14866 1828 14907 1862
rect 14807 1790 14907 1828
rect 14807 1756 14832 1790
rect 14866 1756 14907 1790
rect 14807 1718 14907 1756
rect 14807 1684 14832 1718
rect 14866 1684 14907 1718
rect 14807 1646 14907 1684
rect 14807 1612 14832 1646
rect 14866 1612 14907 1646
rect 14807 1574 14907 1612
rect 14807 1540 14832 1574
rect 14866 1540 14907 1574
rect 14807 1502 14907 1540
rect 14807 1468 14832 1502
rect 14866 1468 14907 1502
rect 14807 1429 14907 1468
rect 14807 1395 14832 1429
rect 14866 1395 14907 1429
rect 14807 1356 14907 1395
rect 14807 1322 14832 1356
rect 14866 1322 14907 1356
rect 14807 1283 14907 1322
rect 14807 1249 14832 1283
rect 14866 1249 14907 1283
rect 14807 1210 14907 1249
rect 14807 1176 14832 1210
rect 14866 1176 14907 1210
rect 14807 1137 14907 1176
rect 14807 1103 14832 1137
rect 14866 1103 14907 1137
rect 14807 1064 14907 1103
rect 14807 1030 14832 1064
rect 14866 1030 14907 1064
rect 14807 991 14907 1030
rect 14807 957 14832 991
rect 14866 957 14907 991
rect 14807 918 14907 957
rect 14807 884 14832 918
rect 14866 884 14907 918
tri 14170 845 14184 859 se
rect 14184 845 14618 859
tri 14793 845 14807 859 se
rect 14807 845 14907 884
rect 303 829 366 845
rect 229 820 366 829
tri 366 820 391 845 sw
rect 517 832 965 845
tri 965 832 978 845 sw
tri 14157 832 14170 845 se
rect 14170 832 14618 845
rect 517 820 14618 832
rect 229 818 391 820
tri 391 818 393 820 sw
rect 517 818 709 820
rect 229 789 393 818
rect 229 755 269 789
rect 303 786 393 789
tri 393 786 425 818 sw
tri 517 786 549 818 ne
rect 549 786 709 818
rect 743 786 782 820
rect 816 786 855 820
rect 889 786 928 820
rect 303 755 425 786
rect 229 748 425 755
tri 425 748 463 786 sw
tri 549 748 587 786 ne
rect 587 748 928 786
rect 229 715 463 748
rect 229 681 269 715
rect 303 714 463 715
tri 463 714 497 748 sw
tri 587 714 621 748 ne
rect 621 714 709 748
rect 743 714 782 748
rect 816 714 855 748
rect 889 714 928 748
rect 14426 818 14618 820
rect 14426 811 14611 818
tri 14611 811 14618 818 nw
tri 14759 811 14793 845 se
rect 14793 811 14832 845
rect 14866 811 14907 845
rect 14426 772 14572 811
tri 14572 772 14611 811 nw
tri 14720 772 14759 811 se
rect 14759 772 14907 811
rect 14426 738 14538 772
tri 14538 738 14572 772 nw
tri 14686 738 14720 772 se
rect 14720 738 14832 772
rect 14866 738 14907 772
rect 14426 714 14502 738
rect 303 702 497 714
tri 497 702 509 714 sw
tri 621 702 633 714 ne
rect 633 702 14502 714
tri 14502 702 14538 738 nw
tri 14650 702 14686 738 se
rect 14686 702 14907 738
rect 303 699 509 702
tri 509 699 512 702 sw
tri 14647 699 14650 702 se
rect 14650 699 14907 702
rect 303 681 512 699
rect 229 665 512 681
tri 512 665 546 699 sw
tri 14613 665 14647 699 se
rect 14647 665 14832 699
rect 14866 665 14907 699
rect 229 641 546 665
rect 229 607 269 641
rect 303 626 546 641
tri 546 626 585 665 sw
tri 14574 626 14613 665 se
rect 14613 626 14907 665
rect 303 607 585 626
rect 229 592 585 607
tri 585 592 619 626 sw
tri 14540 592 14574 626 se
rect 14574 592 14832 626
rect 14866 592 14907 626
rect 229 567 619 592
rect 229 533 269 567
rect 303 553 619 567
tri 619 553 658 592 sw
tri 14501 553 14540 592 se
rect 14540 553 14907 592
rect 303 533 658 553
rect 229 519 658 533
tri 658 519 692 553 sw
tri 14467 519 14501 553 se
rect 14501 519 14832 553
rect 14866 519 14907 553
rect 229 505 692 519
tri 692 505 706 519 sw
tri 14453 505 14467 519 se
rect 14467 505 14907 519
rect 229 497 706 505
rect 229 463 343 497
rect 377 463 419 497
rect 453 463 495 497
rect 529 463 571 497
rect 605 463 648 497
rect 682 481 706 497
tri 706 481 730 505 sw
tri 14435 487 14453 505 se
rect 14453 487 14907 505
tri 14429 481 14435 487 se
rect 14435 481 14907 487
rect 682 463 730 481
rect 229 447 730 463
tri 730 447 764 481 sw
tri 14395 447 14429 481 se
rect 14429 447 14465 481
rect 14499 447 14539 481
rect 14573 447 14613 481
rect 14647 447 14686 481
rect 14720 447 14759 481
rect 14793 447 14907 481
rect 229 402 764 447
tri 764 402 809 447 sw
tri 14389 441 14395 447 se
rect 14395 441 14907 447
tri 14350 402 14389 441 se
rect 14389 402 14907 441
rect 229 375 14907 402
rect 229 341 361 375
rect 395 341 434 375
rect 468 341 507 375
rect 541 341 580 375
rect 614 341 653 375
rect 687 341 726 375
rect 760 341 799 375
rect 833 341 872 375
rect 906 341 945 375
rect 979 341 1018 375
rect 1052 341 1091 375
rect 1125 341 1164 375
rect 1198 341 1237 375
rect 1271 341 1310 375
rect 1344 341 1383 375
rect 1417 341 1456 375
rect 1490 341 1529 375
rect 1563 341 1602 375
rect 1636 341 1675 375
rect 1709 341 1748 375
rect 1782 341 1821 375
rect 1855 341 1894 375
rect 1928 341 1967 375
rect 2001 341 2040 375
rect 2074 341 2113 375
rect 2147 341 2186 375
rect 2220 341 2259 375
rect 2293 341 2332 375
rect 2366 341 2405 375
rect 2439 341 2478 375
rect 2512 341 2551 375
rect 2585 341 2624 375
rect 2658 341 2697 375
rect 2731 341 2770 375
rect 2804 341 2843 375
rect 2877 341 2916 375
rect 2950 341 2989 375
rect 3023 341 3062 375
rect 3096 341 3135 375
rect 3169 341 3208 375
rect 3242 341 3281 375
rect 3315 341 3354 375
rect 3388 341 3427 375
rect 3461 341 3500 375
rect 3534 341 3573 375
rect 3607 341 3646 375
rect 3680 341 3719 375
rect 3753 341 3792 375
rect 3826 341 3865 375
rect 3899 341 3938 375
rect 3972 341 4011 375
rect 4045 341 4084 375
rect 4118 341 4157 375
rect 4191 341 4229 375
rect 4263 341 4301 375
rect 4335 341 4373 375
rect 4407 341 4445 375
rect 4479 341 4517 375
rect 4551 341 4589 375
rect 4623 341 4661 375
rect 4695 341 4733 375
rect 4767 341 4805 375
rect 4839 341 4877 375
rect 4911 341 4949 375
rect 4983 341 5021 375
rect 5055 341 5093 375
rect 5127 341 5165 375
rect 5199 341 5237 375
rect 5271 341 5309 375
rect 5343 341 5381 375
rect 5415 341 5453 375
rect 5487 341 5525 375
rect 5559 341 5597 375
rect 5631 341 5669 375
rect 5703 341 5741 375
rect 5775 341 5813 375
rect 5847 341 5885 375
rect 5919 341 5957 375
rect 5991 341 6029 375
rect 6063 341 6101 375
rect 6135 341 6173 375
rect 6207 341 6245 375
rect 6279 341 6317 375
rect 6351 341 6389 375
rect 6423 341 6461 375
rect 6495 341 6533 375
rect 6567 341 6605 375
rect 6639 341 6677 375
rect 6711 341 6749 375
rect 6783 341 6821 375
rect 6855 341 6893 375
rect 6927 341 6965 375
rect 6999 341 7037 375
rect 7071 341 7109 375
rect 7143 341 7181 375
rect 7215 341 7253 375
rect 7287 341 7325 375
rect 7359 341 7397 375
rect 7431 341 7469 375
rect 7503 341 7541 375
rect 7575 341 7613 375
rect 7647 341 7685 375
rect 7719 341 7757 375
rect 7791 341 7829 375
rect 7863 341 7901 375
rect 7935 341 7973 375
rect 8007 341 8045 375
rect 8079 341 8117 375
rect 8151 341 8189 375
rect 8223 341 8261 375
rect 8295 341 8333 375
rect 8367 341 8405 375
rect 8439 341 8477 375
rect 8511 341 8549 375
rect 8583 341 8621 375
rect 8655 341 8693 375
rect 8727 341 8765 375
rect 8799 341 8837 375
rect 8871 341 8909 375
rect 8943 341 8981 375
rect 9015 341 9053 375
rect 9087 341 9125 375
rect 9159 341 9197 375
rect 9231 341 9269 375
rect 9303 341 9341 375
rect 9375 341 9413 375
rect 9447 341 9485 375
rect 9519 341 9557 375
rect 9591 341 9629 375
rect 9663 341 9701 375
rect 9735 341 9773 375
rect 9807 341 9845 375
rect 9879 341 9917 375
rect 9951 341 9989 375
rect 10023 341 10061 375
rect 10095 341 10133 375
rect 10167 341 10205 375
rect 10239 341 10277 375
rect 10311 341 10349 375
rect 10383 341 10421 375
rect 10455 341 10493 375
rect 10527 341 10565 375
rect 10599 341 10637 375
rect 10671 341 10709 375
rect 10743 341 10781 375
rect 10815 341 10853 375
rect 10887 341 10925 375
rect 10959 341 10997 375
rect 11031 341 11069 375
rect 11103 341 11141 375
rect 11175 341 11213 375
rect 11247 341 11285 375
rect 11319 341 11357 375
rect 11391 341 11429 375
rect 11463 341 11501 375
rect 11535 341 11573 375
rect 11607 341 11645 375
rect 11679 341 11717 375
rect 11751 341 11789 375
rect 11823 341 11861 375
rect 11895 341 11933 375
rect 11967 341 12005 375
rect 12039 341 12077 375
rect 12111 341 12149 375
rect 12183 341 12221 375
rect 12255 341 12293 375
rect 12327 341 12365 375
rect 12399 341 12437 375
rect 12471 341 12509 375
rect 12543 341 12581 375
rect 12615 341 12653 375
rect 12687 341 12725 375
rect 12759 341 12797 375
rect 12831 341 12869 375
rect 12903 341 12941 375
rect 12975 341 13013 375
rect 13047 341 13085 375
rect 13119 341 13157 375
rect 13191 341 13229 375
rect 13263 341 13301 375
rect 13335 341 13373 375
rect 13407 341 13445 375
rect 13479 341 13517 375
rect 13551 341 13589 375
rect 13623 341 13661 375
rect 13695 341 13733 375
rect 13767 341 13805 375
rect 13839 341 13877 375
rect 13911 341 13949 375
rect 13983 341 14021 375
rect 14055 341 14093 375
rect 14127 341 14165 375
rect 14199 341 14237 375
rect 14271 341 14309 375
rect 14343 341 14381 375
rect 14415 341 14453 375
rect 14487 341 14525 375
rect 14559 341 14597 375
rect 14631 341 14669 375
rect 14703 341 14741 375
rect 14775 348 14907 375
rect 15085 348 15097 5062
rect 14775 341 15097 348
rect 229 331 15097 341
rect 39 314 15097 331
<< via1 >>
rect 558 2650 563 2657
rect 563 2650 601 2657
rect 601 2650 610 2657
rect 558 2610 610 2650
rect 558 2605 563 2610
rect 563 2605 601 2610
rect 601 2605 610 2610
rect 646 2605 674 2657
rect 674 2605 698 2657
rect 734 2605 780 2657
rect 780 2605 786 2657
rect 558 2576 563 2592
rect 563 2576 601 2592
rect 601 2576 610 2592
rect 558 2540 610 2576
rect 646 2540 674 2592
rect 674 2540 698 2592
rect 734 2540 780 2592
rect 780 2540 786 2592
rect 558 2502 563 2527
rect 563 2502 601 2527
rect 601 2502 610 2527
rect 558 2475 610 2502
rect 646 2475 674 2527
rect 674 2475 698 2527
rect 734 2475 780 2527
rect 780 2475 786 2527
rect 558 2428 563 2462
rect 563 2428 601 2462
rect 601 2428 610 2462
rect 558 2410 610 2428
rect 646 2410 674 2462
rect 674 2410 698 2462
rect 734 2410 780 2462
rect 780 2410 786 2462
rect 558 2389 610 2397
rect 558 2355 563 2389
rect 563 2355 601 2389
rect 601 2355 610 2389
rect 558 2345 610 2355
rect 646 2345 674 2397
rect 674 2345 698 2397
rect 734 2345 780 2397
rect 780 2345 786 2397
rect 558 2316 610 2332
rect 558 2282 563 2316
rect 563 2282 601 2316
rect 601 2282 610 2316
rect 558 2280 610 2282
rect 646 2280 674 2332
rect 674 2280 698 2332
rect 734 2280 780 2332
rect 780 2280 786 2332
rect 558 2243 610 2267
rect 558 2215 563 2243
rect 563 2215 601 2243
rect 601 2215 610 2243
rect 646 2215 674 2267
rect 674 2215 698 2267
rect 734 2215 780 2267
rect 780 2215 786 2267
rect 558 2170 610 2202
rect 558 2150 563 2170
rect 563 2150 601 2170
rect 601 2150 610 2170
rect 646 2150 674 2202
rect 674 2150 698 2202
rect 734 2150 780 2202
rect 780 2150 786 2202
rect 558 2136 563 2137
rect 563 2136 601 2137
rect 601 2136 610 2137
rect 558 2097 610 2136
rect 558 2085 563 2097
rect 563 2085 601 2097
rect 601 2085 610 2097
rect 646 2085 674 2137
rect 674 2085 698 2137
rect 734 2085 780 2137
rect 780 2085 786 2137
rect 558 2063 563 2072
rect 563 2063 601 2072
rect 601 2063 610 2072
rect 558 2024 610 2063
rect 558 2020 563 2024
rect 563 2020 601 2024
rect 601 2020 610 2024
rect 646 2020 674 2072
rect 674 2020 698 2072
rect 734 2020 780 2072
rect 780 2020 786 2072
rect 558 1990 563 2007
rect 563 1990 601 2007
rect 601 1990 610 2007
rect 558 1955 610 1990
rect 646 1955 674 2007
rect 674 1955 698 2007
rect 734 1955 780 2007
rect 780 1955 786 2007
rect 558 1917 563 1942
rect 563 1917 601 1942
rect 601 1917 610 1942
rect 558 1890 610 1917
rect 646 1890 674 1942
rect 674 1890 698 1942
rect 734 1890 780 1942
rect 780 1890 786 1942
rect 558 1844 563 1877
rect 563 1844 601 1877
rect 601 1844 610 1877
rect 558 1825 610 1844
rect 646 1825 674 1877
rect 674 1825 698 1877
rect 734 1825 780 1877
rect 780 1825 786 1877
rect 558 1805 610 1812
rect 558 1771 563 1805
rect 563 1771 601 1805
rect 601 1771 610 1805
rect 558 1760 610 1771
rect 646 1760 674 1812
rect 674 1760 698 1812
rect 734 1760 780 1812
rect 780 1760 786 1812
rect 558 1732 610 1748
rect 558 1698 563 1732
rect 563 1698 601 1732
rect 601 1698 610 1732
rect 558 1696 610 1698
rect 646 1696 674 1748
rect 674 1696 698 1748
rect 734 1696 780 1748
rect 780 1696 786 1748
rect 558 1659 610 1684
rect 558 1632 563 1659
rect 563 1632 601 1659
rect 601 1632 610 1659
rect 646 1632 674 1684
rect 674 1632 698 1684
rect 734 1632 780 1684
rect 780 1632 786 1684
rect 558 1586 610 1620
rect 558 1568 563 1586
rect 563 1568 601 1586
rect 601 1568 610 1586
rect 646 1568 674 1620
rect 674 1568 698 1620
rect 734 1568 780 1620
rect 780 1568 786 1620
rect 1066 4098 1118 4119
rect 1066 4067 1067 4098
rect 1067 4067 1101 4098
rect 1101 4067 1118 4098
rect 1130 4098 1182 4119
rect 1130 4067 1139 4098
rect 1139 4067 1173 4098
rect 1173 4067 1182 4098
rect 1194 4098 1246 4119
rect 1194 4067 1211 4098
rect 1211 4067 1245 4098
rect 1245 4067 1246 4098
rect 1066 4025 1118 4054
rect 1066 4002 1067 4025
rect 1067 4002 1101 4025
rect 1101 4002 1118 4025
rect 1130 4025 1182 4054
rect 1130 4002 1139 4025
rect 1139 4002 1173 4025
rect 1173 4002 1182 4025
rect 1194 4025 1246 4054
rect 1194 4002 1211 4025
rect 1211 4002 1245 4025
rect 1245 4002 1246 4025
rect 1066 3952 1118 3989
rect 1066 3937 1067 3952
rect 1067 3937 1101 3952
rect 1101 3937 1118 3952
rect 1130 3952 1182 3989
rect 1130 3937 1139 3952
rect 1139 3937 1173 3952
rect 1173 3937 1182 3952
rect 1194 3952 1246 3989
rect 1194 3937 1211 3952
rect 1211 3937 1245 3952
rect 1245 3937 1246 3952
rect 1066 3918 1067 3924
rect 1067 3918 1101 3924
rect 1101 3918 1118 3924
rect 1066 3879 1118 3918
rect 1066 3872 1067 3879
rect 1067 3872 1101 3879
rect 1101 3872 1118 3879
rect 1130 3918 1139 3924
rect 1139 3918 1173 3924
rect 1173 3918 1182 3924
rect 1130 3879 1182 3918
rect 1130 3872 1139 3879
rect 1139 3872 1173 3879
rect 1173 3872 1182 3879
rect 1194 3918 1211 3924
rect 1211 3918 1245 3924
rect 1245 3918 1246 3924
rect 1194 3879 1246 3918
rect 1194 3872 1211 3879
rect 1211 3872 1245 3879
rect 1245 3872 1246 3879
rect 1066 3845 1067 3859
rect 1067 3845 1101 3859
rect 1101 3845 1118 3859
rect 1066 3807 1118 3845
rect 1130 3845 1139 3859
rect 1139 3845 1173 3859
rect 1173 3845 1182 3859
rect 1130 3807 1182 3845
rect 1194 3845 1211 3859
rect 1211 3845 1245 3859
rect 1245 3845 1246 3859
rect 1194 3807 1246 3845
rect 1066 3772 1067 3794
rect 1067 3772 1101 3794
rect 1101 3772 1118 3794
rect 1066 3742 1118 3772
rect 1130 3772 1139 3794
rect 1139 3772 1173 3794
rect 1173 3772 1182 3794
rect 1130 3742 1182 3772
rect 1194 3772 1211 3794
rect 1211 3772 1245 3794
rect 1245 3772 1246 3794
rect 1194 3742 1246 3772
rect 1066 3699 1067 3729
rect 1067 3699 1101 3729
rect 1101 3699 1118 3729
rect 1066 3677 1118 3699
rect 1130 3699 1139 3729
rect 1139 3699 1173 3729
rect 1173 3699 1182 3729
rect 1130 3677 1182 3699
rect 1194 3699 1211 3729
rect 1211 3699 1245 3729
rect 1245 3699 1246 3729
rect 1194 3677 1246 3699
rect 1066 3660 1246 3664
rect 1066 3626 1067 3660
rect 1067 3626 1101 3660
rect 1101 3626 1139 3660
rect 1139 3626 1173 3660
rect 1173 3626 1211 3660
rect 1211 3626 1245 3660
rect 1245 3626 1246 3660
rect 1066 3587 1246 3626
rect 1066 3553 1067 3587
rect 1067 3553 1101 3587
rect 1101 3553 1139 3587
rect 1139 3553 1173 3587
rect 1173 3553 1211 3587
rect 1211 3553 1245 3587
rect 1245 3553 1246 3587
rect 1066 3514 1246 3553
rect 1066 3480 1067 3514
rect 1067 3480 1101 3514
rect 1101 3480 1139 3514
rect 1139 3480 1173 3514
rect 1173 3480 1211 3514
rect 1211 3480 1245 3514
rect 1245 3480 1246 3514
rect 1066 3441 1246 3480
rect 1066 3407 1067 3441
rect 1067 3407 1101 3441
rect 1101 3407 1139 3441
rect 1139 3407 1173 3441
rect 1173 3407 1211 3441
rect 1211 3407 1245 3441
rect 1245 3407 1246 3441
rect 1066 3368 1246 3407
rect 1066 3334 1067 3368
rect 1067 3334 1101 3368
rect 1101 3334 1139 3368
rect 1139 3334 1173 3368
rect 1173 3334 1211 3368
rect 1211 3334 1245 3368
rect 1245 3334 1246 3368
rect 1066 3295 1246 3334
rect 1066 3261 1067 3295
rect 1067 3261 1101 3295
rect 1101 3261 1139 3295
rect 1139 3261 1173 3295
rect 1173 3261 1211 3295
rect 1211 3261 1245 3295
rect 1245 3261 1246 3295
rect 1066 3222 1246 3261
rect 1066 3188 1067 3222
rect 1067 3188 1101 3222
rect 1101 3188 1139 3222
rect 1139 3188 1173 3222
rect 1173 3188 1211 3222
rect 1211 3188 1245 3222
rect 1245 3188 1246 3222
rect 1066 3149 1246 3188
rect 1066 3115 1067 3149
rect 1067 3115 1101 3149
rect 1101 3115 1139 3149
rect 1139 3115 1173 3149
rect 1173 3115 1211 3149
rect 1211 3115 1245 3149
rect 1245 3115 1246 3149
rect 1066 3076 1246 3115
rect 1066 3042 1067 3076
rect 1067 3042 1101 3076
rect 1101 3042 1139 3076
rect 1139 3042 1173 3076
rect 1173 3042 1211 3076
rect 1211 3042 1245 3076
rect 1245 3042 1246 3076
rect 1066 3003 1246 3042
rect 1066 2972 1067 3003
rect 1067 2972 1101 3003
rect 1101 2972 1139 3003
rect 1139 2972 1173 3003
rect 1173 2972 1211 3003
rect 1211 2972 1245 3003
rect 1245 2972 1246 3003
rect 1562 2628 1614 2657
rect 1562 2605 1563 2628
rect 1563 2605 1597 2628
rect 1597 2605 1614 2628
rect 1626 2628 1678 2657
rect 1626 2605 1635 2628
rect 1635 2605 1669 2628
rect 1669 2605 1678 2628
rect 1690 2628 1742 2657
rect 1690 2605 1707 2628
rect 1707 2605 1741 2628
rect 1741 2605 1742 2628
rect 1562 2540 1614 2592
rect 1626 2556 1678 2592
rect 1626 2540 1635 2556
rect 1635 2540 1669 2556
rect 1669 2540 1678 2556
rect 1690 2540 1742 2592
rect 1562 2518 1614 2527
rect 1626 2522 1635 2527
rect 1635 2522 1669 2527
rect 1669 2522 1678 2527
rect 1626 2518 1678 2522
rect 1690 2518 1742 2527
rect 1562 2475 1563 2518
rect 1563 2475 1614 2518
rect 1626 2475 1678 2518
rect 1690 2475 1741 2518
rect 1741 2475 1742 2518
rect 1562 2410 1563 2462
rect 1563 2410 1614 2462
rect 1626 2410 1678 2462
rect 1690 2410 1741 2462
rect 1741 2410 1742 2462
rect 1562 2345 1563 2397
rect 1563 2345 1614 2397
rect 1626 2345 1678 2397
rect 1690 2345 1741 2397
rect 1741 2345 1742 2397
rect 1562 2280 1563 2332
rect 1563 2280 1614 2332
rect 1626 2280 1678 2332
rect 1690 2280 1741 2332
rect 1741 2280 1742 2332
rect 1562 2215 1563 2267
rect 1563 2215 1614 2267
rect 1626 2215 1678 2267
rect 1690 2215 1741 2267
rect 1741 2215 1742 2267
rect 1562 2150 1563 2202
rect 1563 2150 1614 2202
rect 1626 2150 1678 2202
rect 1690 2150 1741 2202
rect 1741 2150 1742 2202
rect 1562 2085 1563 2137
rect 1563 2085 1614 2137
rect 1626 2085 1678 2137
rect 1690 2085 1741 2137
rect 1741 2085 1742 2137
rect 1562 2020 1563 2072
rect 1563 2020 1614 2072
rect 1626 2020 1678 2072
rect 1690 2020 1741 2072
rect 1741 2020 1742 2072
rect 1562 1955 1563 2007
rect 1563 1955 1614 2007
rect 1626 1955 1678 2007
rect 1690 1955 1741 2007
rect 1741 1955 1742 2007
rect 1562 1890 1563 1942
rect 1563 1890 1614 1942
rect 1626 1890 1678 1942
rect 1690 1890 1741 1942
rect 1741 1890 1742 1942
rect 1562 1825 1563 1877
rect 1563 1825 1614 1877
rect 1626 1825 1678 1877
rect 1690 1825 1741 1877
rect 1741 1825 1742 1877
rect 1562 1620 1563 1812
rect 1563 1620 1741 1812
rect 1741 1620 1742 1812
rect 1562 1586 1635 1620
rect 1635 1586 1669 1620
rect 1669 1586 1742 1620
rect 1562 1568 1742 1586
rect 2058 4098 2110 4119
rect 2058 4067 2059 4098
rect 2059 4067 2093 4098
rect 2093 4067 2110 4098
rect 2122 4098 2174 4119
rect 2122 4067 2131 4098
rect 2131 4067 2165 4098
rect 2165 4067 2174 4098
rect 2186 4098 2238 4119
rect 2186 4067 2203 4098
rect 2203 4067 2237 4098
rect 2237 4067 2238 4098
rect 2058 4025 2110 4054
rect 2058 4002 2059 4025
rect 2059 4002 2093 4025
rect 2093 4002 2110 4025
rect 2122 4025 2174 4054
rect 2122 4002 2131 4025
rect 2131 4002 2165 4025
rect 2165 4002 2174 4025
rect 2186 4025 2238 4054
rect 2186 4002 2203 4025
rect 2203 4002 2237 4025
rect 2237 4002 2238 4025
rect 2058 3952 2110 3989
rect 2058 3937 2059 3952
rect 2059 3937 2093 3952
rect 2093 3937 2110 3952
rect 2122 3952 2174 3989
rect 2122 3937 2131 3952
rect 2131 3937 2165 3952
rect 2165 3937 2174 3952
rect 2186 3952 2238 3989
rect 2186 3937 2203 3952
rect 2203 3937 2237 3952
rect 2237 3937 2238 3952
rect 2058 3918 2059 3924
rect 2059 3918 2093 3924
rect 2093 3918 2110 3924
rect 2058 3879 2110 3918
rect 2058 3872 2059 3879
rect 2059 3872 2093 3879
rect 2093 3872 2110 3879
rect 2122 3918 2131 3924
rect 2131 3918 2165 3924
rect 2165 3918 2174 3924
rect 2122 3879 2174 3918
rect 2122 3872 2131 3879
rect 2131 3872 2165 3879
rect 2165 3872 2174 3879
rect 2186 3918 2203 3924
rect 2203 3918 2237 3924
rect 2237 3918 2238 3924
rect 2186 3879 2238 3918
rect 2186 3872 2203 3879
rect 2203 3872 2237 3879
rect 2237 3872 2238 3879
rect 2058 3845 2059 3859
rect 2059 3845 2093 3859
rect 2093 3845 2110 3859
rect 2058 3807 2110 3845
rect 2122 3845 2131 3859
rect 2131 3845 2165 3859
rect 2165 3845 2174 3859
rect 2122 3807 2174 3845
rect 2186 3845 2203 3859
rect 2203 3845 2237 3859
rect 2237 3845 2238 3859
rect 2186 3807 2238 3845
rect 2058 3772 2059 3794
rect 2059 3772 2093 3794
rect 2093 3772 2110 3794
rect 2058 3742 2110 3772
rect 2122 3772 2131 3794
rect 2131 3772 2165 3794
rect 2165 3772 2174 3794
rect 2122 3742 2174 3772
rect 2186 3772 2203 3794
rect 2203 3772 2237 3794
rect 2237 3772 2238 3794
rect 2186 3742 2238 3772
rect 2058 3699 2059 3729
rect 2059 3699 2093 3729
rect 2093 3699 2110 3729
rect 2058 3677 2110 3699
rect 2122 3699 2131 3729
rect 2131 3699 2165 3729
rect 2165 3699 2174 3729
rect 2122 3677 2174 3699
rect 2186 3699 2203 3729
rect 2203 3699 2237 3729
rect 2237 3699 2238 3729
rect 2186 3677 2238 3699
rect 2058 3660 2238 3664
rect 2058 3626 2059 3660
rect 2059 3626 2093 3660
rect 2093 3626 2131 3660
rect 2131 3626 2165 3660
rect 2165 3626 2203 3660
rect 2203 3626 2237 3660
rect 2237 3626 2238 3660
rect 2058 3587 2238 3626
rect 2058 3553 2059 3587
rect 2059 3553 2093 3587
rect 2093 3553 2131 3587
rect 2131 3553 2165 3587
rect 2165 3553 2203 3587
rect 2203 3553 2237 3587
rect 2237 3553 2238 3587
rect 2058 3514 2238 3553
rect 2058 3480 2059 3514
rect 2059 3480 2093 3514
rect 2093 3480 2131 3514
rect 2131 3480 2165 3514
rect 2165 3480 2203 3514
rect 2203 3480 2237 3514
rect 2237 3480 2238 3514
rect 2058 3441 2238 3480
rect 2058 3407 2059 3441
rect 2059 3407 2093 3441
rect 2093 3407 2131 3441
rect 2131 3407 2165 3441
rect 2165 3407 2203 3441
rect 2203 3407 2237 3441
rect 2237 3407 2238 3441
rect 2058 3368 2238 3407
rect 2058 3334 2059 3368
rect 2059 3334 2093 3368
rect 2093 3334 2131 3368
rect 2131 3334 2165 3368
rect 2165 3334 2203 3368
rect 2203 3334 2237 3368
rect 2237 3334 2238 3368
rect 2058 3295 2238 3334
rect 2058 3261 2059 3295
rect 2059 3261 2093 3295
rect 2093 3261 2131 3295
rect 2131 3261 2165 3295
rect 2165 3261 2203 3295
rect 2203 3261 2237 3295
rect 2237 3261 2238 3295
rect 2058 3222 2238 3261
rect 2058 3188 2059 3222
rect 2059 3188 2093 3222
rect 2093 3188 2131 3222
rect 2131 3188 2165 3222
rect 2165 3188 2203 3222
rect 2203 3188 2237 3222
rect 2237 3188 2238 3222
rect 2058 3149 2238 3188
rect 2058 3115 2059 3149
rect 2059 3115 2093 3149
rect 2093 3115 2131 3149
rect 2131 3115 2165 3149
rect 2165 3115 2203 3149
rect 2203 3115 2237 3149
rect 2237 3115 2238 3149
rect 2058 3076 2238 3115
rect 2058 3042 2059 3076
rect 2059 3042 2093 3076
rect 2093 3042 2131 3076
rect 2131 3042 2165 3076
rect 2165 3042 2203 3076
rect 2203 3042 2237 3076
rect 2237 3042 2238 3076
rect 2058 3003 2238 3042
rect 2058 2972 2059 3003
rect 2059 2972 2093 3003
rect 2093 2972 2131 3003
rect 2131 2972 2165 3003
rect 2165 2972 2203 3003
rect 2203 2972 2237 3003
rect 2237 2972 2238 3003
rect 2554 2628 2606 2657
rect 2554 2605 2555 2628
rect 2555 2605 2589 2628
rect 2589 2605 2606 2628
rect 2618 2628 2670 2657
rect 2618 2605 2627 2628
rect 2627 2605 2661 2628
rect 2661 2605 2670 2628
rect 2682 2628 2734 2657
rect 2682 2605 2699 2628
rect 2699 2605 2733 2628
rect 2733 2605 2734 2628
rect 2554 2540 2606 2592
rect 2618 2556 2670 2592
rect 2618 2540 2627 2556
rect 2627 2540 2661 2556
rect 2661 2540 2670 2556
rect 2682 2540 2734 2592
rect 2554 2518 2606 2527
rect 2618 2522 2627 2527
rect 2627 2522 2661 2527
rect 2661 2522 2670 2527
rect 2618 2518 2670 2522
rect 2682 2518 2734 2527
rect 2554 2475 2555 2518
rect 2555 2475 2606 2518
rect 2618 2475 2670 2518
rect 2682 2475 2733 2518
rect 2733 2475 2734 2518
rect 2554 2410 2555 2462
rect 2555 2410 2606 2462
rect 2618 2410 2670 2462
rect 2682 2410 2733 2462
rect 2733 2410 2734 2462
rect 2554 2345 2555 2397
rect 2555 2345 2606 2397
rect 2618 2345 2670 2397
rect 2682 2345 2733 2397
rect 2733 2345 2734 2397
rect 2554 2280 2555 2332
rect 2555 2280 2606 2332
rect 2618 2280 2670 2332
rect 2682 2280 2733 2332
rect 2733 2280 2734 2332
rect 2554 2215 2555 2267
rect 2555 2215 2606 2267
rect 2618 2215 2670 2267
rect 2682 2215 2733 2267
rect 2733 2215 2734 2267
rect 2554 2150 2555 2202
rect 2555 2150 2606 2202
rect 2618 2150 2670 2202
rect 2682 2150 2733 2202
rect 2733 2150 2734 2202
rect 2554 2085 2555 2137
rect 2555 2085 2606 2137
rect 2618 2085 2670 2137
rect 2682 2085 2733 2137
rect 2733 2085 2734 2137
rect 2554 2020 2555 2072
rect 2555 2020 2606 2072
rect 2618 2020 2670 2072
rect 2682 2020 2733 2072
rect 2733 2020 2734 2072
rect 2554 1955 2555 2007
rect 2555 1955 2606 2007
rect 2618 1955 2670 2007
rect 2682 1955 2733 2007
rect 2733 1955 2734 2007
rect 2554 1890 2555 1942
rect 2555 1890 2606 1942
rect 2618 1890 2670 1942
rect 2682 1890 2733 1942
rect 2733 1890 2734 1942
rect 2554 1825 2555 1877
rect 2555 1825 2606 1877
rect 2618 1825 2670 1877
rect 2682 1825 2733 1877
rect 2733 1825 2734 1877
rect 2554 1620 2555 1812
rect 2555 1620 2733 1812
rect 2733 1620 2734 1812
rect 2554 1586 2627 1620
rect 2627 1586 2661 1620
rect 2661 1586 2734 1620
rect 2554 1568 2734 1586
rect 3050 4098 3102 4119
rect 3050 4067 3051 4098
rect 3051 4067 3085 4098
rect 3085 4067 3102 4098
rect 3114 4098 3166 4119
rect 3114 4067 3123 4098
rect 3123 4067 3157 4098
rect 3157 4067 3166 4098
rect 3178 4098 3230 4119
rect 3178 4067 3195 4098
rect 3195 4067 3229 4098
rect 3229 4067 3230 4098
rect 3050 4025 3102 4054
rect 3050 4002 3051 4025
rect 3051 4002 3085 4025
rect 3085 4002 3102 4025
rect 3114 4025 3166 4054
rect 3114 4002 3123 4025
rect 3123 4002 3157 4025
rect 3157 4002 3166 4025
rect 3178 4025 3230 4054
rect 3178 4002 3195 4025
rect 3195 4002 3229 4025
rect 3229 4002 3230 4025
rect 3050 3952 3102 3989
rect 3050 3937 3051 3952
rect 3051 3937 3085 3952
rect 3085 3937 3102 3952
rect 3114 3952 3166 3989
rect 3114 3937 3123 3952
rect 3123 3937 3157 3952
rect 3157 3937 3166 3952
rect 3178 3952 3230 3989
rect 3178 3937 3195 3952
rect 3195 3937 3229 3952
rect 3229 3937 3230 3952
rect 3050 3918 3051 3924
rect 3051 3918 3085 3924
rect 3085 3918 3102 3924
rect 3050 3879 3102 3918
rect 3050 3872 3051 3879
rect 3051 3872 3085 3879
rect 3085 3872 3102 3879
rect 3114 3918 3123 3924
rect 3123 3918 3157 3924
rect 3157 3918 3166 3924
rect 3114 3879 3166 3918
rect 3114 3872 3123 3879
rect 3123 3872 3157 3879
rect 3157 3872 3166 3879
rect 3178 3918 3195 3924
rect 3195 3918 3229 3924
rect 3229 3918 3230 3924
rect 3178 3879 3230 3918
rect 3178 3872 3195 3879
rect 3195 3872 3229 3879
rect 3229 3872 3230 3879
rect 3050 3845 3051 3859
rect 3051 3845 3085 3859
rect 3085 3845 3102 3859
rect 3050 3807 3102 3845
rect 3114 3845 3123 3859
rect 3123 3845 3157 3859
rect 3157 3845 3166 3859
rect 3114 3807 3166 3845
rect 3178 3845 3195 3859
rect 3195 3845 3229 3859
rect 3229 3845 3230 3859
rect 3178 3807 3230 3845
rect 3050 3772 3051 3794
rect 3051 3772 3085 3794
rect 3085 3772 3102 3794
rect 3050 3742 3102 3772
rect 3114 3772 3123 3794
rect 3123 3772 3157 3794
rect 3157 3772 3166 3794
rect 3114 3742 3166 3772
rect 3178 3772 3195 3794
rect 3195 3772 3229 3794
rect 3229 3772 3230 3794
rect 3178 3742 3230 3772
rect 3050 3699 3051 3729
rect 3051 3699 3085 3729
rect 3085 3699 3102 3729
rect 3050 3677 3102 3699
rect 3114 3699 3123 3729
rect 3123 3699 3157 3729
rect 3157 3699 3166 3729
rect 3114 3677 3166 3699
rect 3178 3699 3195 3729
rect 3195 3699 3229 3729
rect 3229 3699 3230 3729
rect 3178 3677 3230 3699
rect 3050 3660 3230 3664
rect 3050 3626 3051 3660
rect 3051 3626 3085 3660
rect 3085 3626 3123 3660
rect 3123 3626 3157 3660
rect 3157 3626 3195 3660
rect 3195 3626 3229 3660
rect 3229 3626 3230 3660
rect 3050 3587 3230 3626
rect 3050 3553 3051 3587
rect 3051 3553 3085 3587
rect 3085 3553 3123 3587
rect 3123 3553 3157 3587
rect 3157 3553 3195 3587
rect 3195 3553 3229 3587
rect 3229 3553 3230 3587
rect 3050 3514 3230 3553
rect 3050 3480 3051 3514
rect 3051 3480 3085 3514
rect 3085 3480 3123 3514
rect 3123 3480 3157 3514
rect 3157 3480 3195 3514
rect 3195 3480 3229 3514
rect 3229 3480 3230 3514
rect 3050 3441 3230 3480
rect 3050 3407 3051 3441
rect 3051 3407 3085 3441
rect 3085 3407 3123 3441
rect 3123 3407 3157 3441
rect 3157 3407 3195 3441
rect 3195 3407 3229 3441
rect 3229 3407 3230 3441
rect 3050 3368 3230 3407
rect 3050 3334 3051 3368
rect 3051 3334 3085 3368
rect 3085 3334 3123 3368
rect 3123 3334 3157 3368
rect 3157 3334 3195 3368
rect 3195 3334 3229 3368
rect 3229 3334 3230 3368
rect 3050 3295 3230 3334
rect 3050 3261 3051 3295
rect 3051 3261 3085 3295
rect 3085 3261 3123 3295
rect 3123 3261 3157 3295
rect 3157 3261 3195 3295
rect 3195 3261 3229 3295
rect 3229 3261 3230 3295
rect 3050 3222 3230 3261
rect 3050 3188 3051 3222
rect 3051 3188 3085 3222
rect 3085 3188 3123 3222
rect 3123 3188 3157 3222
rect 3157 3188 3195 3222
rect 3195 3188 3229 3222
rect 3229 3188 3230 3222
rect 3050 3149 3230 3188
rect 3050 3115 3051 3149
rect 3051 3115 3085 3149
rect 3085 3115 3123 3149
rect 3123 3115 3157 3149
rect 3157 3115 3195 3149
rect 3195 3115 3229 3149
rect 3229 3115 3230 3149
rect 3050 3076 3230 3115
rect 3050 3042 3051 3076
rect 3051 3042 3085 3076
rect 3085 3042 3123 3076
rect 3123 3042 3157 3076
rect 3157 3042 3195 3076
rect 3195 3042 3229 3076
rect 3229 3042 3230 3076
rect 3050 3003 3230 3042
rect 3050 2972 3051 3003
rect 3051 2972 3085 3003
rect 3085 2972 3123 3003
rect 3123 2972 3157 3003
rect 3157 2972 3195 3003
rect 3195 2972 3229 3003
rect 3229 2972 3230 3003
rect 3546 2628 3598 2657
rect 3546 2605 3547 2628
rect 3547 2605 3581 2628
rect 3581 2605 3598 2628
rect 3610 2628 3662 2657
rect 3610 2605 3619 2628
rect 3619 2605 3653 2628
rect 3653 2605 3662 2628
rect 3674 2628 3726 2657
rect 3674 2605 3691 2628
rect 3691 2605 3725 2628
rect 3725 2605 3726 2628
rect 3546 2540 3598 2592
rect 3610 2556 3662 2592
rect 3610 2540 3619 2556
rect 3619 2540 3653 2556
rect 3653 2540 3662 2556
rect 3674 2540 3726 2592
rect 3546 2518 3598 2527
rect 3610 2522 3619 2527
rect 3619 2522 3653 2527
rect 3653 2522 3662 2527
rect 3610 2518 3662 2522
rect 3674 2518 3726 2527
rect 3546 2475 3547 2518
rect 3547 2475 3598 2518
rect 3610 2475 3662 2518
rect 3674 2475 3725 2518
rect 3725 2475 3726 2518
rect 3546 2410 3547 2462
rect 3547 2410 3598 2462
rect 3610 2410 3662 2462
rect 3674 2410 3725 2462
rect 3725 2410 3726 2462
rect 3546 2345 3547 2397
rect 3547 2345 3598 2397
rect 3610 2345 3662 2397
rect 3674 2345 3725 2397
rect 3725 2345 3726 2397
rect 3546 2280 3547 2332
rect 3547 2280 3598 2332
rect 3610 2280 3662 2332
rect 3674 2280 3725 2332
rect 3725 2280 3726 2332
rect 3546 2215 3547 2267
rect 3547 2215 3598 2267
rect 3610 2215 3662 2267
rect 3674 2215 3725 2267
rect 3725 2215 3726 2267
rect 3546 2150 3547 2202
rect 3547 2150 3598 2202
rect 3610 2150 3662 2202
rect 3674 2150 3725 2202
rect 3725 2150 3726 2202
rect 3546 2085 3547 2137
rect 3547 2085 3598 2137
rect 3610 2085 3662 2137
rect 3674 2085 3725 2137
rect 3725 2085 3726 2137
rect 3546 2020 3547 2072
rect 3547 2020 3598 2072
rect 3610 2020 3662 2072
rect 3674 2020 3725 2072
rect 3725 2020 3726 2072
rect 3546 1955 3547 2007
rect 3547 1955 3598 2007
rect 3610 1955 3662 2007
rect 3674 1955 3725 2007
rect 3725 1955 3726 2007
rect 3546 1890 3547 1942
rect 3547 1890 3598 1942
rect 3610 1890 3662 1942
rect 3674 1890 3725 1942
rect 3725 1890 3726 1942
rect 3546 1825 3547 1877
rect 3547 1825 3598 1877
rect 3610 1825 3662 1877
rect 3674 1825 3725 1877
rect 3725 1825 3726 1877
rect 3546 1620 3547 1812
rect 3547 1620 3725 1812
rect 3725 1620 3726 1812
rect 3546 1586 3619 1620
rect 3619 1586 3653 1620
rect 3653 1586 3726 1620
rect 3546 1568 3726 1586
rect 4042 4098 4094 4119
rect 4042 4067 4043 4098
rect 4043 4067 4077 4098
rect 4077 4067 4094 4098
rect 4106 4098 4158 4119
rect 4106 4067 4115 4098
rect 4115 4067 4149 4098
rect 4149 4067 4158 4098
rect 4170 4098 4222 4119
rect 4170 4067 4187 4098
rect 4187 4067 4221 4098
rect 4221 4067 4222 4098
rect 4042 4025 4094 4054
rect 4042 4002 4043 4025
rect 4043 4002 4077 4025
rect 4077 4002 4094 4025
rect 4106 4025 4158 4054
rect 4106 4002 4115 4025
rect 4115 4002 4149 4025
rect 4149 4002 4158 4025
rect 4170 4025 4222 4054
rect 4170 4002 4187 4025
rect 4187 4002 4221 4025
rect 4221 4002 4222 4025
rect 4042 3952 4094 3989
rect 4042 3937 4043 3952
rect 4043 3937 4077 3952
rect 4077 3937 4094 3952
rect 4106 3952 4158 3989
rect 4106 3937 4115 3952
rect 4115 3937 4149 3952
rect 4149 3937 4158 3952
rect 4170 3952 4222 3989
rect 4170 3937 4187 3952
rect 4187 3937 4221 3952
rect 4221 3937 4222 3952
rect 4042 3918 4043 3924
rect 4043 3918 4077 3924
rect 4077 3918 4094 3924
rect 4042 3879 4094 3918
rect 4042 3872 4043 3879
rect 4043 3872 4077 3879
rect 4077 3872 4094 3879
rect 4106 3918 4115 3924
rect 4115 3918 4149 3924
rect 4149 3918 4158 3924
rect 4106 3879 4158 3918
rect 4106 3872 4115 3879
rect 4115 3872 4149 3879
rect 4149 3872 4158 3879
rect 4170 3918 4187 3924
rect 4187 3918 4221 3924
rect 4221 3918 4222 3924
rect 4170 3879 4222 3918
rect 4170 3872 4187 3879
rect 4187 3872 4221 3879
rect 4221 3872 4222 3879
rect 4042 3845 4043 3859
rect 4043 3845 4077 3859
rect 4077 3845 4094 3859
rect 4042 3807 4094 3845
rect 4106 3845 4115 3859
rect 4115 3845 4149 3859
rect 4149 3845 4158 3859
rect 4106 3807 4158 3845
rect 4170 3845 4187 3859
rect 4187 3845 4221 3859
rect 4221 3845 4222 3859
rect 4170 3807 4222 3845
rect 4042 3772 4043 3794
rect 4043 3772 4077 3794
rect 4077 3772 4094 3794
rect 4042 3742 4094 3772
rect 4106 3772 4115 3794
rect 4115 3772 4149 3794
rect 4149 3772 4158 3794
rect 4106 3742 4158 3772
rect 4170 3772 4187 3794
rect 4187 3772 4221 3794
rect 4221 3772 4222 3794
rect 4170 3742 4222 3772
rect 4042 3699 4043 3729
rect 4043 3699 4077 3729
rect 4077 3699 4094 3729
rect 4042 3677 4094 3699
rect 4106 3699 4115 3729
rect 4115 3699 4149 3729
rect 4149 3699 4158 3729
rect 4106 3677 4158 3699
rect 4170 3699 4187 3729
rect 4187 3699 4221 3729
rect 4221 3699 4222 3729
rect 4170 3677 4222 3699
rect 4042 3660 4222 3664
rect 4042 3626 4043 3660
rect 4043 3626 4077 3660
rect 4077 3626 4115 3660
rect 4115 3626 4149 3660
rect 4149 3626 4187 3660
rect 4187 3626 4221 3660
rect 4221 3626 4222 3660
rect 4042 3587 4222 3626
rect 4042 3553 4043 3587
rect 4043 3553 4077 3587
rect 4077 3553 4115 3587
rect 4115 3553 4149 3587
rect 4149 3553 4187 3587
rect 4187 3553 4221 3587
rect 4221 3553 4222 3587
rect 4042 3514 4222 3553
rect 4042 3480 4043 3514
rect 4043 3480 4077 3514
rect 4077 3480 4115 3514
rect 4115 3480 4149 3514
rect 4149 3480 4187 3514
rect 4187 3480 4221 3514
rect 4221 3480 4222 3514
rect 4042 3441 4222 3480
rect 4042 3407 4043 3441
rect 4043 3407 4077 3441
rect 4077 3407 4115 3441
rect 4115 3407 4149 3441
rect 4149 3407 4187 3441
rect 4187 3407 4221 3441
rect 4221 3407 4222 3441
rect 4042 3368 4222 3407
rect 4042 3334 4043 3368
rect 4043 3334 4077 3368
rect 4077 3334 4115 3368
rect 4115 3334 4149 3368
rect 4149 3334 4187 3368
rect 4187 3334 4221 3368
rect 4221 3334 4222 3368
rect 4042 3295 4222 3334
rect 4042 3261 4043 3295
rect 4043 3261 4077 3295
rect 4077 3261 4115 3295
rect 4115 3261 4149 3295
rect 4149 3261 4187 3295
rect 4187 3261 4221 3295
rect 4221 3261 4222 3295
rect 4042 3222 4222 3261
rect 4042 3188 4043 3222
rect 4043 3188 4077 3222
rect 4077 3188 4115 3222
rect 4115 3188 4149 3222
rect 4149 3188 4187 3222
rect 4187 3188 4221 3222
rect 4221 3188 4222 3222
rect 4042 3149 4222 3188
rect 4042 3115 4043 3149
rect 4043 3115 4077 3149
rect 4077 3115 4115 3149
rect 4115 3115 4149 3149
rect 4149 3115 4187 3149
rect 4187 3115 4221 3149
rect 4221 3115 4222 3149
rect 4042 3076 4222 3115
rect 4042 3042 4043 3076
rect 4043 3042 4077 3076
rect 4077 3042 4115 3076
rect 4115 3042 4149 3076
rect 4149 3042 4187 3076
rect 4187 3042 4221 3076
rect 4221 3042 4222 3076
rect 4042 3003 4222 3042
rect 4042 2972 4043 3003
rect 4043 2972 4077 3003
rect 4077 2972 4115 3003
rect 4115 2972 4149 3003
rect 4149 2972 4187 3003
rect 4187 2972 4221 3003
rect 4221 2972 4222 3003
rect 4538 2628 4590 2657
rect 4538 2605 4539 2628
rect 4539 2605 4573 2628
rect 4573 2605 4590 2628
rect 4602 2628 4654 2657
rect 4602 2605 4611 2628
rect 4611 2605 4645 2628
rect 4645 2605 4654 2628
rect 4666 2628 4718 2657
rect 4666 2605 4683 2628
rect 4683 2605 4717 2628
rect 4717 2605 4718 2628
rect 4538 2540 4590 2592
rect 4602 2556 4654 2592
rect 4602 2540 4611 2556
rect 4611 2540 4645 2556
rect 4645 2540 4654 2556
rect 4666 2540 4718 2592
rect 4538 2518 4590 2527
rect 4602 2522 4611 2527
rect 4611 2522 4645 2527
rect 4645 2522 4654 2527
rect 4602 2518 4654 2522
rect 4666 2518 4718 2527
rect 4538 2475 4539 2518
rect 4539 2475 4590 2518
rect 4602 2475 4654 2518
rect 4666 2475 4717 2518
rect 4717 2475 4718 2518
rect 4538 2410 4539 2462
rect 4539 2410 4590 2462
rect 4602 2410 4654 2462
rect 4666 2410 4717 2462
rect 4717 2410 4718 2462
rect 4538 2345 4539 2397
rect 4539 2345 4590 2397
rect 4602 2345 4654 2397
rect 4666 2345 4717 2397
rect 4717 2345 4718 2397
rect 4538 2280 4539 2332
rect 4539 2280 4590 2332
rect 4602 2280 4654 2332
rect 4666 2280 4717 2332
rect 4717 2280 4718 2332
rect 4538 2215 4539 2267
rect 4539 2215 4590 2267
rect 4602 2215 4654 2267
rect 4666 2215 4717 2267
rect 4717 2215 4718 2267
rect 4538 2150 4539 2202
rect 4539 2150 4590 2202
rect 4602 2150 4654 2202
rect 4666 2150 4717 2202
rect 4717 2150 4718 2202
rect 4538 2085 4539 2137
rect 4539 2085 4590 2137
rect 4602 2085 4654 2137
rect 4666 2085 4717 2137
rect 4717 2085 4718 2137
rect 4538 2020 4539 2072
rect 4539 2020 4590 2072
rect 4602 2020 4654 2072
rect 4666 2020 4717 2072
rect 4717 2020 4718 2072
rect 4538 1955 4539 2007
rect 4539 1955 4590 2007
rect 4602 1955 4654 2007
rect 4666 1955 4717 2007
rect 4717 1955 4718 2007
rect 4538 1890 4539 1942
rect 4539 1890 4590 1942
rect 4602 1890 4654 1942
rect 4666 1890 4717 1942
rect 4717 1890 4718 1942
rect 4538 1825 4539 1877
rect 4539 1825 4590 1877
rect 4602 1825 4654 1877
rect 4666 1825 4717 1877
rect 4717 1825 4718 1877
rect 4538 1620 4539 1812
rect 4539 1620 4717 1812
rect 4717 1620 4718 1812
rect 4538 1586 4611 1620
rect 4611 1586 4645 1620
rect 4645 1586 4718 1620
rect 4538 1568 4718 1586
rect 5034 4098 5086 4119
rect 5034 4067 5035 4098
rect 5035 4067 5069 4098
rect 5069 4067 5086 4098
rect 5098 4098 5150 4119
rect 5098 4067 5107 4098
rect 5107 4067 5141 4098
rect 5141 4067 5150 4098
rect 5162 4098 5214 4119
rect 5162 4067 5179 4098
rect 5179 4067 5213 4098
rect 5213 4067 5214 4098
rect 5034 4025 5086 4054
rect 5034 4002 5035 4025
rect 5035 4002 5069 4025
rect 5069 4002 5086 4025
rect 5098 4025 5150 4054
rect 5098 4002 5107 4025
rect 5107 4002 5141 4025
rect 5141 4002 5150 4025
rect 5162 4025 5214 4054
rect 5162 4002 5179 4025
rect 5179 4002 5213 4025
rect 5213 4002 5214 4025
rect 5034 3952 5086 3989
rect 5034 3937 5035 3952
rect 5035 3937 5069 3952
rect 5069 3937 5086 3952
rect 5098 3952 5150 3989
rect 5098 3937 5107 3952
rect 5107 3937 5141 3952
rect 5141 3937 5150 3952
rect 5162 3952 5214 3989
rect 5162 3937 5179 3952
rect 5179 3937 5213 3952
rect 5213 3937 5214 3952
rect 5034 3918 5035 3924
rect 5035 3918 5069 3924
rect 5069 3918 5086 3924
rect 5034 3879 5086 3918
rect 5034 3872 5035 3879
rect 5035 3872 5069 3879
rect 5069 3872 5086 3879
rect 5098 3918 5107 3924
rect 5107 3918 5141 3924
rect 5141 3918 5150 3924
rect 5098 3879 5150 3918
rect 5098 3872 5107 3879
rect 5107 3872 5141 3879
rect 5141 3872 5150 3879
rect 5162 3918 5179 3924
rect 5179 3918 5213 3924
rect 5213 3918 5214 3924
rect 5162 3879 5214 3918
rect 5162 3872 5179 3879
rect 5179 3872 5213 3879
rect 5213 3872 5214 3879
rect 5034 3845 5035 3859
rect 5035 3845 5069 3859
rect 5069 3845 5086 3859
rect 5034 3807 5086 3845
rect 5098 3845 5107 3859
rect 5107 3845 5141 3859
rect 5141 3845 5150 3859
rect 5098 3807 5150 3845
rect 5162 3845 5179 3859
rect 5179 3845 5213 3859
rect 5213 3845 5214 3859
rect 5162 3807 5214 3845
rect 5034 3772 5035 3794
rect 5035 3772 5069 3794
rect 5069 3772 5086 3794
rect 5034 3742 5086 3772
rect 5098 3772 5107 3794
rect 5107 3772 5141 3794
rect 5141 3772 5150 3794
rect 5098 3742 5150 3772
rect 5162 3772 5179 3794
rect 5179 3772 5213 3794
rect 5213 3772 5214 3794
rect 5162 3742 5214 3772
rect 5034 3699 5035 3729
rect 5035 3699 5069 3729
rect 5069 3699 5086 3729
rect 5034 3677 5086 3699
rect 5098 3699 5107 3729
rect 5107 3699 5141 3729
rect 5141 3699 5150 3729
rect 5098 3677 5150 3699
rect 5162 3699 5179 3729
rect 5179 3699 5213 3729
rect 5213 3699 5214 3729
rect 5162 3677 5214 3699
rect 5034 3660 5214 3664
rect 5034 3626 5035 3660
rect 5035 3626 5069 3660
rect 5069 3626 5107 3660
rect 5107 3626 5141 3660
rect 5141 3626 5179 3660
rect 5179 3626 5213 3660
rect 5213 3626 5214 3660
rect 5034 3587 5214 3626
rect 5034 3553 5035 3587
rect 5035 3553 5069 3587
rect 5069 3553 5107 3587
rect 5107 3553 5141 3587
rect 5141 3553 5179 3587
rect 5179 3553 5213 3587
rect 5213 3553 5214 3587
rect 5034 3514 5214 3553
rect 5034 3480 5035 3514
rect 5035 3480 5069 3514
rect 5069 3480 5107 3514
rect 5107 3480 5141 3514
rect 5141 3480 5179 3514
rect 5179 3480 5213 3514
rect 5213 3480 5214 3514
rect 5034 3441 5214 3480
rect 5034 3407 5035 3441
rect 5035 3407 5069 3441
rect 5069 3407 5107 3441
rect 5107 3407 5141 3441
rect 5141 3407 5179 3441
rect 5179 3407 5213 3441
rect 5213 3407 5214 3441
rect 5034 3368 5214 3407
rect 5034 3334 5035 3368
rect 5035 3334 5069 3368
rect 5069 3334 5107 3368
rect 5107 3334 5141 3368
rect 5141 3334 5179 3368
rect 5179 3334 5213 3368
rect 5213 3334 5214 3368
rect 5034 3295 5214 3334
rect 5034 3261 5035 3295
rect 5035 3261 5069 3295
rect 5069 3261 5107 3295
rect 5107 3261 5141 3295
rect 5141 3261 5179 3295
rect 5179 3261 5213 3295
rect 5213 3261 5214 3295
rect 5034 3222 5214 3261
rect 5034 3188 5035 3222
rect 5035 3188 5069 3222
rect 5069 3188 5107 3222
rect 5107 3188 5141 3222
rect 5141 3188 5179 3222
rect 5179 3188 5213 3222
rect 5213 3188 5214 3222
rect 5034 3149 5214 3188
rect 5034 3115 5035 3149
rect 5035 3115 5069 3149
rect 5069 3115 5107 3149
rect 5107 3115 5141 3149
rect 5141 3115 5179 3149
rect 5179 3115 5213 3149
rect 5213 3115 5214 3149
rect 5034 3076 5214 3115
rect 5034 3042 5035 3076
rect 5035 3042 5069 3076
rect 5069 3042 5107 3076
rect 5107 3042 5141 3076
rect 5141 3042 5179 3076
rect 5179 3042 5213 3076
rect 5213 3042 5214 3076
rect 5034 3003 5214 3042
rect 5034 2972 5035 3003
rect 5035 2972 5069 3003
rect 5069 2972 5107 3003
rect 5107 2972 5141 3003
rect 5141 2972 5179 3003
rect 5179 2972 5213 3003
rect 5213 2972 5214 3003
rect 5530 2628 5582 2657
rect 5530 2605 5531 2628
rect 5531 2605 5565 2628
rect 5565 2605 5582 2628
rect 5594 2628 5646 2657
rect 5594 2605 5603 2628
rect 5603 2605 5637 2628
rect 5637 2605 5646 2628
rect 5658 2628 5710 2657
rect 5658 2605 5675 2628
rect 5675 2605 5709 2628
rect 5709 2605 5710 2628
rect 5530 2540 5582 2592
rect 5594 2556 5646 2592
rect 5594 2540 5603 2556
rect 5603 2540 5637 2556
rect 5637 2540 5646 2556
rect 5658 2540 5710 2592
rect 5530 2518 5582 2527
rect 5594 2522 5603 2527
rect 5603 2522 5637 2527
rect 5637 2522 5646 2527
rect 5594 2518 5646 2522
rect 5658 2518 5710 2527
rect 5530 2475 5531 2518
rect 5531 2475 5582 2518
rect 5594 2475 5646 2518
rect 5658 2475 5709 2518
rect 5709 2475 5710 2518
rect 5530 2410 5531 2462
rect 5531 2410 5582 2462
rect 5594 2410 5646 2462
rect 5658 2410 5709 2462
rect 5709 2410 5710 2462
rect 5530 2345 5531 2397
rect 5531 2345 5582 2397
rect 5594 2345 5646 2397
rect 5658 2345 5709 2397
rect 5709 2345 5710 2397
rect 5530 2280 5531 2332
rect 5531 2280 5582 2332
rect 5594 2280 5646 2332
rect 5658 2280 5709 2332
rect 5709 2280 5710 2332
rect 5530 2215 5531 2267
rect 5531 2215 5582 2267
rect 5594 2215 5646 2267
rect 5658 2215 5709 2267
rect 5709 2215 5710 2267
rect 5530 2150 5531 2202
rect 5531 2150 5582 2202
rect 5594 2150 5646 2202
rect 5658 2150 5709 2202
rect 5709 2150 5710 2202
rect 5530 2085 5531 2137
rect 5531 2085 5582 2137
rect 5594 2085 5646 2137
rect 5658 2085 5709 2137
rect 5709 2085 5710 2137
rect 5530 2020 5531 2072
rect 5531 2020 5582 2072
rect 5594 2020 5646 2072
rect 5658 2020 5709 2072
rect 5709 2020 5710 2072
rect 5530 1955 5531 2007
rect 5531 1955 5582 2007
rect 5594 1955 5646 2007
rect 5658 1955 5709 2007
rect 5709 1955 5710 2007
rect 5530 1890 5531 1942
rect 5531 1890 5582 1942
rect 5594 1890 5646 1942
rect 5658 1890 5709 1942
rect 5709 1890 5710 1942
rect 5530 1825 5531 1877
rect 5531 1825 5582 1877
rect 5594 1825 5646 1877
rect 5658 1825 5709 1877
rect 5709 1825 5710 1877
rect 5530 1620 5531 1812
rect 5531 1620 5709 1812
rect 5709 1620 5710 1812
rect 5530 1586 5603 1620
rect 5603 1586 5637 1620
rect 5637 1586 5710 1620
rect 5530 1568 5710 1586
rect 6026 4098 6078 4119
rect 6026 4067 6027 4098
rect 6027 4067 6061 4098
rect 6061 4067 6078 4098
rect 6090 4098 6142 4119
rect 6090 4067 6099 4098
rect 6099 4067 6133 4098
rect 6133 4067 6142 4098
rect 6154 4098 6206 4119
rect 6154 4067 6171 4098
rect 6171 4067 6205 4098
rect 6205 4067 6206 4098
rect 6026 4025 6078 4054
rect 6026 4002 6027 4025
rect 6027 4002 6061 4025
rect 6061 4002 6078 4025
rect 6090 4025 6142 4054
rect 6090 4002 6099 4025
rect 6099 4002 6133 4025
rect 6133 4002 6142 4025
rect 6154 4025 6206 4054
rect 6154 4002 6171 4025
rect 6171 4002 6205 4025
rect 6205 4002 6206 4025
rect 6026 3952 6078 3989
rect 6026 3937 6027 3952
rect 6027 3937 6061 3952
rect 6061 3937 6078 3952
rect 6090 3952 6142 3989
rect 6090 3937 6099 3952
rect 6099 3937 6133 3952
rect 6133 3937 6142 3952
rect 6154 3952 6206 3989
rect 6154 3937 6171 3952
rect 6171 3937 6205 3952
rect 6205 3937 6206 3952
rect 6026 3918 6027 3924
rect 6027 3918 6061 3924
rect 6061 3918 6078 3924
rect 6026 3879 6078 3918
rect 6026 3872 6027 3879
rect 6027 3872 6061 3879
rect 6061 3872 6078 3879
rect 6090 3918 6099 3924
rect 6099 3918 6133 3924
rect 6133 3918 6142 3924
rect 6090 3879 6142 3918
rect 6090 3872 6099 3879
rect 6099 3872 6133 3879
rect 6133 3872 6142 3879
rect 6154 3918 6171 3924
rect 6171 3918 6205 3924
rect 6205 3918 6206 3924
rect 6154 3879 6206 3918
rect 6154 3872 6171 3879
rect 6171 3872 6205 3879
rect 6205 3872 6206 3879
rect 6026 3845 6027 3859
rect 6027 3845 6061 3859
rect 6061 3845 6078 3859
rect 6026 3807 6078 3845
rect 6090 3845 6099 3859
rect 6099 3845 6133 3859
rect 6133 3845 6142 3859
rect 6090 3807 6142 3845
rect 6154 3845 6171 3859
rect 6171 3845 6205 3859
rect 6205 3845 6206 3859
rect 6154 3807 6206 3845
rect 6026 3772 6027 3794
rect 6027 3772 6061 3794
rect 6061 3772 6078 3794
rect 6026 3742 6078 3772
rect 6090 3772 6099 3794
rect 6099 3772 6133 3794
rect 6133 3772 6142 3794
rect 6090 3742 6142 3772
rect 6154 3772 6171 3794
rect 6171 3772 6205 3794
rect 6205 3772 6206 3794
rect 6154 3742 6206 3772
rect 6026 3699 6027 3729
rect 6027 3699 6061 3729
rect 6061 3699 6078 3729
rect 6026 3677 6078 3699
rect 6090 3699 6099 3729
rect 6099 3699 6133 3729
rect 6133 3699 6142 3729
rect 6090 3677 6142 3699
rect 6154 3699 6171 3729
rect 6171 3699 6205 3729
rect 6205 3699 6206 3729
rect 6154 3677 6206 3699
rect 6026 3660 6206 3664
rect 6026 3626 6027 3660
rect 6027 3626 6061 3660
rect 6061 3626 6099 3660
rect 6099 3626 6133 3660
rect 6133 3626 6171 3660
rect 6171 3626 6205 3660
rect 6205 3626 6206 3660
rect 6026 3587 6206 3626
rect 6026 3553 6027 3587
rect 6027 3553 6061 3587
rect 6061 3553 6099 3587
rect 6099 3553 6133 3587
rect 6133 3553 6171 3587
rect 6171 3553 6205 3587
rect 6205 3553 6206 3587
rect 6026 3514 6206 3553
rect 6026 3480 6027 3514
rect 6027 3480 6061 3514
rect 6061 3480 6099 3514
rect 6099 3480 6133 3514
rect 6133 3480 6171 3514
rect 6171 3480 6205 3514
rect 6205 3480 6206 3514
rect 6026 3441 6206 3480
rect 6026 3407 6027 3441
rect 6027 3407 6061 3441
rect 6061 3407 6099 3441
rect 6099 3407 6133 3441
rect 6133 3407 6171 3441
rect 6171 3407 6205 3441
rect 6205 3407 6206 3441
rect 6026 3368 6206 3407
rect 6026 3334 6027 3368
rect 6027 3334 6061 3368
rect 6061 3334 6099 3368
rect 6099 3334 6133 3368
rect 6133 3334 6171 3368
rect 6171 3334 6205 3368
rect 6205 3334 6206 3368
rect 6026 3295 6206 3334
rect 6026 3261 6027 3295
rect 6027 3261 6061 3295
rect 6061 3261 6099 3295
rect 6099 3261 6133 3295
rect 6133 3261 6171 3295
rect 6171 3261 6205 3295
rect 6205 3261 6206 3295
rect 6026 3222 6206 3261
rect 6026 3188 6027 3222
rect 6027 3188 6061 3222
rect 6061 3188 6099 3222
rect 6099 3188 6133 3222
rect 6133 3188 6171 3222
rect 6171 3188 6205 3222
rect 6205 3188 6206 3222
rect 6026 3149 6206 3188
rect 6026 3115 6027 3149
rect 6027 3115 6061 3149
rect 6061 3115 6099 3149
rect 6099 3115 6133 3149
rect 6133 3115 6171 3149
rect 6171 3115 6205 3149
rect 6205 3115 6206 3149
rect 6026 3076 6206 3115
rect 6026 3042 6027 3076
rect 6027 3042 6061 3076
rect 6061 3042 6099 3076
rect 6099 3042 6133 3076
rect 6133 3042 6171 3076
rect 6171 3042 6205 3076
rect 6205 3042 6206 3076
rect 6026 3003 6206 3042
rect 6026 2972 6027 3003
rect 6027 2972 6061 3003
rect 6061 2972 6099 3003
rect 6099 2972 6133 3003
rect 6133 2972 6171 3003
rect 6171 2972 6205 3003
rect 6205 2972 6206 3003
rect 6522 2628 6574 2657
rect 6522 2605 6523 2628
rect 6523 2605 6557 2628
rect 6557 2605 6574 2628
rect 6586 2628 6638 2657
rect 6586 2605 6595 2628
rect 6595 2605 6629 2628
rect 6629 2605 6638 2628
rect 6650 2628 6702 2657
rect 6650 2605 6667 2628
rect 6667 2605 6701 2628
rect 6701 2605 6702 2628
rect 6522 2540 6574 2592
rect 6586 2556 6638 2592
rect 6586 2540 6595 2556
rect 6595 2540 6629 2556
rect 6629 2540 6638 2556
rect 6650 2540 6702 2592
rect 6522 2518 6574 2527
rect 6586 2522 6595 2527
rect 6595 2522 6629 2527
rect 6629 2522 6638 2527
rect 6586 2518 6638 2522
rect 6650 2518 6702 2527
rect 6522 2475 6523 2518
rect 6523 2475 6574 2518
rect 6586 2475 6638 2518
rect 6650 2475 6701 2518
rect 6701 2475 6702 2518
rect 6522 2410 6523 2462
rect 6523 2410 6574 2462
rect 6586 2410 6638 2462
rect 6650 2410 6701 2462
rect 6701 2410 6702 2462
rect 6522 2345 6523 2397
rect 6523 2345 6574 2397
rect 6586 2345 6638 2397
rect 6650 2345 6701 2397
rect 6701 2345 6702 2397
rect 6522 2280 6523 2332
rect 6523 2280 6574 2332
rect 6586 2280 6638 2332
rect 6650 2280 6701 2332
rect 6701 2280 6702 2332
rect 6522 2215 6523 2267
rect 6523 2215 6574 2267
rect 6586 2215 6638 2267
rect 6650 2215 6701 2267
rect 6701 2215 6702 2267
rect 6522 2150 6523 2202
rect 6523 2150 6574 2202
rect 6586 2150 6638 2202
rect 6650 2150 6701 2202
rect 6701 2150 6702 2202
rect 6522 2085 6523 2137
rect 6523 2085 6574 2137
rect 6586 2085 6638 2137
rect 6650 2085 6701 2137
rect 6701 2085 6702 2137
rect 6522 2020 6523 2072
rect 6523 2020 6574 2072
rect 6586 2020 6638 2072
rect 6650 2020 6701 2072
rect 6701 2020 6702 2072
rect 6522 1955 6523 2007
rect 6523 1955 6574 2007
rect 6586 1955 6638 2007
rect 6650 1955 6701 2007
rect 6701 1955 6702 2007
rect 6522 1890 6523 1942
rect 6523 1890 6574 1942
rect 6586 1890 6638 1942
rect 6650 1890 6701 1942
rect 6701 1890 6702 1942
rect 6522 1825 6523 1877
rect 6523 1825 6574 1877
rect 6586 1825 6638 1877
rect 6650 1825 6701 1877
rect 6701 1825 6702 1877
rect 6522 1620 6523 1812
rect 6523 1620 6701 1812
rect 6701 1620 6702 1812
rect 6522 1586 6595 1620
rect 6595 1586 6629 1620
rect 6629 1586 6702 1620
rect 6522 1568 6702 1586
rect 7018 4098 7070 4119
rect 7018 4067 7019 4098
rect 7019 4067 7053 4098
rect 7053 4067 7070 4098
rect 7082 4098 7134 4119
rect 7082 4067 7091 4098
rect 7091 4067 7125 4098
rect 7125 4067 7134 4098
rect 7146 4098 7198 4119
rect 7146 4067 7163 4098
rect 7163 4067 7197 4098
rect 7197 4067 7198 4098
rect 7018 4025 7070 4054
rect 7018 4002 7019 4025
rect 7019 4002 7053 4025
rect 7053 4002 7070 4025
rect 7082 4025 7134 4054
rect 7082 4002 7091 4025
rect 7091 4002 7125 4025
rect 7125 4002 7134 4025
rect 7146 4025 7198 4054
rect 7146 4002 7163 4025
rect 7163 4002 7197 4025
rect 7197 4002 7198 4025
rect 7018 3952 7070 3989
rect 7018 3937 7019 3952
rect 7019 3937 7053 3952
rect 7053 3937 7070 3952
rect 7082 3952 7134 3989
rect 7082 3937 7091 3952
rect 7091 3937 7125 3952
rect 7125 3937 7134 3952
rect 7146 3952 7198 3989
rect 7146 3937 7163 3952
rect 7163 3937 7197 3952
rect 7197 3937 7198 3952
rect 7018 3918 7019 3924
rect 7019 3918 7053 3924
rect 7053 3918 7070 3924
rect 7018 3879 7070 3918
rect 7018 3872 7019 3879
rect 7019 3872 7053 3879
rect 7053 3872 7070 3879
rect 7082 3918 7091 3924
rect 7091 3918 7125 3924
rect 7125 3918 7134 3924
rect 7082 3879 7134 3918
rect 7082 3872 7091 3879
rect 7091 3872 7125 3879
rect 7125 3872 7134 3879
rect 7146 3918 7163 3924
rect 7163 3918 7197 3924
rect 7197 3918 7198 3924
rect 7146 3879 7198 3918
rect 7146 3872 7163 3879
rect 7163 3872 7197 3879
rect 7197 3872 7198 3879
rect 7018 3845 7019 3859
rect 7019 3845 7053 3859
rect 7053 3845 7070 3859
rect 7018 3807 7070 3845
rect 7082 3845 7091 3859
rect 7091 3845 7125 3859
rect 7125 3845 7134 3859
rect 7082 3807 7134 3845
rect 7146 3845 7163 3859
rect 7163 3845 7197 3859
rect 7197 3845 7198 3859
rect 7146 3807 7198 3845
rect 7018 3772 7019 3794
rect 7019 3772 7053 3794
rect 7053 3772 7070 3794
rect 7018 3742 7070 3772
rect 7082 3772 7091 3794
rect 7091 3772 7125 3794
rect 7125 3772 7134 3794
rect 7082 3742 7134 3772
rect 7146 3772 7163 3794
rect 7163 3772 7197 3794
rect 7197 3772 7198 3794
rect 7146 3742 7198 3772
rect 7018 3699 7019 3729
rect 7019 3699 7053 3729
rect 7053 3699 7070 3729
rect 7018 3677 7070 3699
rect 7082 3699 7091 3729
rect 7091 3699 7125 3729
rect 7125 3699 7134 3729
rect 7082 3677 7134 3699
rect 7146 3699 7163 3729
rect 7163 3699 7197 3729
rect 7197 3699 7198 3729
rect 7146 3677 7198 3699
rect 7018 3660 7198 3664
rect 7018 3626 7019 3660
rect 7019 3626 7053 3660
rect 7053 3626 7091 3660
rect 7091 3626 7125 3660
rect 7125 3626 7163 3660
rect 7163 3626 7197 3660
rect 7197 3626 7198 3660
rect 7018 3587 7198 3626
rect 7018 3553 7019 3587
rect 7019 3553 7053 3587
rect 7053 3553 7091 3587
rect 7091 3553 7125 3587
rect 7125 3553 7163 3587
rect 7163 3553 7197 3587
rect 7197 3553 7198 3587
rect 7018 3514 7198 3553
rect 7018 3480 7019 3514
rect 7019 3480 7053 3514
rect 7053 3480 7091 3514
rect 7091 3480 7125 3514
rect 7125 3480 7163 3514
rect 7163 3480 7197 3514
rect 7197 3480 7198 3514
rect 7018 3441 7198 3480
rect 7018 3407 7019 3441
rect 7019 3407 7053 3441
rect 7053 3407 7091 3441
rect 7091 3407 7125 3441
rect 7125 3407 7163 3441
rect 7163 3407 7197 3441
rect 7197 3407 7198 3441
rect 7018 3368 7198 3407
rect 7018 3334 7019 3368
rect 7019 3334 7053 3368
rect 7053 3334 7091 3368
rect 7091 3334 7125 3368
rect 7125 3334 7163 3368
rect 7163 3334 7197 3368
rect 7197 3334 7198 3368
rect 7018 3295 7198 3334
rect 7018 3261 7019 3295
rect 7019 3261 7053 3295
rect 7053 3261 7091 3295
rect 7091 3261 7125 3295
rect 7125 3261 7163 3295
rect 7163 3261 7197 3295
rect 7197 3261 7198 3295
rect 7018 3222 7198 3261
rect 7018 3188 7019 3222
rect 7019 3188 7053 3222
rect 7053 3188 7091 3222
rect 7091 3188 7125 3222
rect 7125 3188 7163 3222
rect 7163 3188 7197 3222
rect 7197 3188 7198 3222
rect 7018 3149 7198 3188
rect 7018 3115 7019 3149
rect 7019 3115 7053 3149
rect 7053 3115 7091 3149
rect 7091 3115 7125 3149
rect 7125 3115 7163 3149
rect 7163 3115 7197 3149
rect 7197 3115 7198 3149
rect 7018 3076 7198 3115
rect 7018 3042 7019 3076
rect 7019 3042 7053 3076
rect 7053 3042 7091 3076
rect 7091 3042 7125 3076
rect 7125 3042 7163 3076
rect 7163 3042 7197 3076
rect 7197 3042 7198 3076
rect 7018 3003 7198 3042
rect 7018 2972 7019 3003
rect 7019 2972 7053 3003
rect 7053 2972 7091 3003
rect 7091 2972 7125 3003
rect 7125 2972 7163 3003
rect 7163 2972 7197 3003
rect 7197 2972 7198 3003
rect 7514 2628 7566 2657
rect 7514 2605 7515 2628
rect 7515 2605 7549 2628
rect 7549 2605 7566 2628
rect 7578 2628 7630 2657
rect 7578 2605 7587 2628
rect 7587 2605 7621 2628
rect 7621 2605 7630 2628
rect 7642 2628 7694 2657
rect 7642 2605 7659 2628
rect 7659 2605 7693 2628
rect 7693 2605 7694 2628
rect 7514 2540 7566 2592
rect 7578 2556 7630 2592
rect 7578 2540 7587 2556
rect 7587 2540 7621 2556
rect 7621 2540 7630 2556
rect 7642 2540 7694 2592
rect 7514 2518 7566 2527
rect 7578 2522 7587 2527
rect 7587 2522 7621 2527
rect 7621 2522 7630 2527
rect 7578 2518 7630 2522
rect 7642 2518 7694 2527
rect 7514 2475 7515 2518
rect 7515 2475 7566 2518
rect 7578 2475 7630 2518
rect 7642 2475 7693 2518
rect 7693 2475 7694 2518
rect 7514 2410 7515 2462
rect 7515 2410 7566 2462
rect 7578 2410 7630 2462
rect 7642 2410 7693 2462
rect 7693 2410 7694 2462
rect 7514 2345 7515 2397
rect 7515 2345 7566 2397
rect 7578 2345 7630 2397
rect 7642 2345 7693 2397
rect 7693 2345 7694 2397
rect 7514 2280 7515 2332
rect 7515 2280 7566 2332
rect 7578 2280 7630 2332
rect 7642 2280 7693 2332
rect 7693 2280 7694 2332
rect 7514 2215 7515 2267
rect 7515 2215 7566 2267
rect 7578 2215 7630 2267
rect 7642 2215 7693 2267
rect 7693 2215 7694 2267
rect 7514 2150 7515 2202
rect 7515 2150 7566 2202
rect 7578 2150 7630 2202
rect 7642 2150 7693 2202
rect 7693 2150 7694 2202
rect 7514 2085 7515 2137
rect 7515 2085 7566 2137
rect 7578 2085 7630 2137
rect 7642 2085 7693 2137
rect 7693 2085 7694 2137
rect 7514 2020 7515 2072
rect 7515 2020 7566 2072
rect 7578 2020 7630 2072
rect 7642 2020 7693 2072
rect 7693 2020 7694 2072
rect 7514 1955 7515 2007
rect 7515 1955 7566 2007
rect 7578 1955 7630 2007
rect 7642 1955 7693 2007
rect 7693 1955 7694 2007
rect 7514 1890 7515 1942
rect 7515 1890 7566 1942
rect 7578 1890 7630 1942
rect 7642 1890 7693 1942
rect 7693 1890 7694 1942
rect 7514 1825 7515 1877
rect 7515 1825 7566 1877
rect 7578 1825 7630 1877
rect 7642 1825 7693 1877
rect 7693 1825 7694 1877
rect 7514 1620 7515 1812
rect 7515 1620 7693 1812
rect 7693 1620 7694 1812
rect 7514 1586 7587 1620
rect 7587 1586 7621 1620
rect 7621 1586 7694 1620
rect 7514 1568 7694 1586
rect 8010 4098 8062 4119
rect 8010 4067 8011 4098
rect 8011 4067 8045 4098
rect 8045 4067 8062 4098
rect 8074 4098 8126 4119
rect 8074 4067 8083 4098
rect 8083 4067 8117 4098
rect 8117 4067 8126 4098
rect 8138 4098 8190 4119
rect 8138 4067 8155 4098
rect 8155 4067 8189 4098
rect 8189 4067 8190 4098
rect 8010 4025 8062 4054
rect 8010 4002 8011 4025
rect 8011 4002 8045 4025
rect 8045 4002 8062 4025
rect 8074 4025 8126 4054
rect 8074 4002 8083 4025
rect 8083 4002 8117 4025
rect 8117 4002 8126 4025
rect 8138 4025 8190 4054
rect 8138 4002 8155 4025
rect 8155 4002 8189 4025
rect 8189 4002 8190 4025
rect 8010 3952 8062 3989
rect 8010 3937 8011 3952
rect 8011 3937 8045 3952
rect 8045 3937 8062 3952
rect 8074 3952 8126 3989
rect 8074 3937 8083 3952
rect 8083 3937 8117 3952
rect 8117 3937 8126 3952
rect 8138 3952 8190 3989
rect 8138 3937 8155 3952
rect 8155 3937 8189 3952
rect 8189 3937 8190 3952
rect 8010 3918 8011 3924
rect 8011 3918 8045 3924
rect 8045 3918 8062 3924
rect 8010 3879 8062 3918
rect 8010 3872 8011 3879
rect 8011 3872 8045 3879
rect 8045 3872 8062 3879
rect 8074 3918 8083 3924
rect 8083 3918 8117 3924
rect 8117 3918 8126 3924
rect 8074 3879 8126 3918
rect 8074 3872 8083 3879
rect 8083 3872 8117 3879
rect 8117 3872 8126 3879
rect 8138 3918 8155 3924
rect 8155 3918 8189 3924
rect 8189 3918 8190 3924
rect 8138 3879 8190 3918
rect 8138 3872 8155 3879
rect 8155 3872 8189 3879
rect 8189 3872 8190 3879
rect 8010 3845 8011 3859
rect 8011 3845 8045 3859
rect 8045 3845 8062 3859
rect 8010 3807 8062 3845
rect 8074 3845 8083 3859
rect 8083 3845 8117 3859
rect 8117 3845 8126 3859
rect 8074 3807 8126 3845
rect 8138 3845 8155 3859
rect 8155 3845 8189 3859
rect 8189 3845 8190 3859
rect 8138 3807 8190 3845
rect 8010 3772 8011 3794
rect 8011 3772 8045 3794
rect 8045 3772 8062 3794
rect 8010 3742 8062 3772
rect 8074 3772 8083 3794
rect 8083 3772 8117 3794
rect 8117 3772 8126 3794
rect 8074 3742 8126 3772
rect 8138 3772 8155 3794
rect 8155 3772 8189 3794
rect 8189 3772 8190 3794
rect 8138 3742 8190 3772
rect 8010 3699 8011 3729
rect 8011 3699 8045 3729
rect 8045 3699 8062 3729
rect 8010 3677 8062 3699
rect 8074 3699 8083 3729
rect 8083 3699 8117 3729
rect 8117 3699 8126 3729
rect 8074 3677 8126 3699
rect 8138 3699 8155 3729
rect 8155 3699 8189 3729
rect 8189 3699 8190 3729
rect 8138 3677 8190 3699
rect 8010 3660 8190 3664
rect 8010 3626 8011 3660
rect 8011 3626 8045 3660
rect 8045 3626 8083 3660
rect 8083 3626 8117 3660
rect 8117 3626 8155 3660
rect 8155 3626 8189 3660
rect 8189 3626 8190 3660
rect 8010 3587 8190 3626
rect 8010 3553 8011 3587
rect 8011 3553 8045 3587
rect 8045 3553 8083 3587
rect 8083 3553 8117 3587
rect 8117 3553 8155 3587
rect 8155 3553 8189 3587
rect 8189 3553 8190 3587
rect 8010 3514 8190 3553
rect 8010 3480 8011 3514
rect 8011 3480 8045 3514
rect 8045 3480 8083 3514
rect 8083 3480 8117 3514
rect 8117 3480 8155 3514
rect 8155 3480 8189 3514
rect 8189 3480 8190 3514
rect 8010 3441 8190 3480
rect 8010 3407 8011 3441
rect 8011 3407 8045 3441
rect 8045 3407 8083 3441
rect 8083 3407 8117 3441
rect 8117 3407 8155 3441
rect 8155 3407 8189 3441
rect 8189 3407 8190 3441
rect 8010 3368 8190 3407
rect 8010 3334 8011 3368
rect 8011 3334 8045 3368
rect 8045 3334 8083 3368
rect 8083 3334 8117 3368
rect 8117 3334 8155 3368
rect 8155 3334 8189 3368
rect 8189 3334 8190 3368
rect 8010 3295 8190 3334
rect 8010 3261 8011 3295
rect 8011 3261 8045 3295
rect 8045 3261 8083 3295
rect 8083 3261 8117 3295
rect 8117 3261 8155 3295
rect 8155 3261 8189 3295
rect 8189 3261 8190 3295
rect 8010 3222 8190 3261
rect 8010 3188 8011 3222
rect 8011 3188 8045 3222
rect 8045 3188 8083 3222
rect 8083 3188 8117 3222
rect 8117 3188 8155 3222
rect 8155 3188 8189 3222
rect 8189 3188 8190 3222
rect 8010 3149 8190 3188
rect 8010 3115 8011 3149
rect 8011 3115 8045 3149
rect 8045 3115 8083 3149
rect 8083 3115 8117 3149
rect 8117 3115 8155 3149
rect 8155 3115 8189 3149
rect 8189 3115 8190 3149
rect 8010 3076 8190 3115
rect 8010 3042 8011 3076
rect 8011 3042 8045 3076
rect 8045 3042 8083 3076
rect 8083 3042 8117 3076
rect 8117 3042 8155 3076
rect 8155 3042 8189 3076
rect 8189 3042 8190 3076
rect 8010 3003 8190 3042
rect 8010 2972 8011 3003
rect 8011 2972 8045 3003
rect 8045 2972 8083 3003
rect 8083 2972 8117 3003
rect 8117 2972 8155 3003
rect 8155 2972 8189 3003
rect 8189 2972 8190 3003
rect 8506 2628 8558 2657
rect 8506 2605 8507 2628
rect 8507 2605 8541 2628
rect 8541 2605 8558 2628
rect 8570 2628 8622 2657
rect 8570 2605 8579 2628
rect 8579 2605 8613 2628
rect 8613 2605 8622 2628
rect 8634 2628 8686 2657
rect 8634 2605 8651 2628
rect 8651 2605 8685 2628
rect 8685 2605 8686 2628
rect 8506 2540 8558 2592
rect 8570 2556 8622 2592
rect 8570 2540 8579 2556
rect 8579 2540 8613 2556
rect 8613 2540 8622 2556
rect 8634 2540 8686 2592
rect 8506 2518 8558 2527
rect 8570 2522 8579 2527
rect 8579 2522 8613 2527
rect 8613 2522 8622 2527
rect 8570 2518 8622 2522
rect 8634 2518 8686 2527
rect 8506 2475 8507 2518
rect 8507 2475 8558 2518
rect 8570 2475 8622 2518
rect 8634 2475 8685 2518
rect 8685 2475 8686 2518
rect 8506 2410 8507 2462
rect 8507 2410 8558 2462
rect 8570 2410 8622 2462
rect 8634 2410 8685 2462
rect 8685 2410 8686 2462
rect 8506 2345 8507 2397
rect 8507 2345 8558 2397
rect 8570 2345 8622 2397
rect 8634 2345 8685 2397
rect 8685 2345 8686 2397
rect 8506 2280 8507 2332
rect 8507 2280 8558 2332
rect 8570 2280 8622 2332
rect 8634 2280 8685 2332
rect 8685 2280 8686 2332
rect 8506 2215 8507 2267
rect 8507 2215 8558 2267
rect 8570 2215 8622 2267
rect 8634 2215 8685 2267
rect 8685 2215 8686 2267
rect 8506 2150 8507 2202
rect 8507 2150 8558 2202
rect 8570 2150 8622 2202
rect 8634 2150 8685 2202
rect 8685 2150 8686 2202
rect 8506 2085 8507 2137
rect 8507 2085 8558 2137
rect 8570 2085 8622 2137
rect 8634 2085 8685 2137
rect 8685 2085 8686 2137
rect 8506 2020 8507 2072
rect 8507 2020 8558 2072
rect 8570 2020 8622 2072
rect 8634 2020 8685 2072
rect 8685 2020 8686 2072
rect 8506 1955 8507 2007
rect 8507 1955 8558 2007
rect 8570 1955 8622 2007
rect 8634 1955 8685 2007
rect 8685 1955 8686 2007
rect 8506 1890 8507 1942
rect 8507 1890 8558 1942
rect 8570 1890 8622 1942
rect 8634 1890 8685 1942
rect 8685 1890 8686 1942
rect 8506 1825 8507 1877
rect 8507 1825 8558 1877
rect 8570 1825 8622 1877
rect 8634 1825 8685 1877
rect 8685 1825 8686 1877
rect 8506 1620 8507 1812
rect 8507 1620 8685 1812
rect 8685 1620 8686 1812
rect 8506 1586 8579 1620
rect 8579 1586 8613 1620
rect 8613 1586 8686 1620
rect 8506 1568 8686 1586
rect 9002 4098 9054 4119
rect 9002 4067 9003 4098
rect 9003 4067 9037 4098
rect 9037 4067 9054 4098
rect 9066 4098 9118 4119
rect 9066 4067 9075 4098
rect 9075 4067 9109 4098
rect 9109 4067 9118 4098
rect 9130 4098 9182 4119
rect 9130 4067 9147 4098
rect 9147 4067 9181 4098
rect 9181 4067 9182 4098
rect 9002 4025 9054 4054
rect 9002 4002 9003 4025
rect 9003 4002 9037 4025
rect 9037 4002 9054 4025
rect 9066 4025 9118 4054
rect 9066 4002 9075 4025
rect 9075 4002 9109 4025
rect 9109 4002 9118 4025
rect 9130 4025 9182 4054
rect 9130 4002 9147 4025
rect 9147 4002 9181 4025
rect 9181 4002 9182 4025
rect 9002 3952 9054 3989
rect 9002 3937 9003 3952
rect 9003 3937 9037 3952
rect 9037 3937 9054 3952
rect 9066 3952 9118 3989
rect 9066 3937 9075 3952
rect 9075 3937 9109 3952
rect 9109 3937 9118 3952
rect 9130 3952 9182 3989
rect 9130 3937 9147 3952
rect 9147 3937 9181 3952
rect 9181 3937 9182 3952
rect 9002 3918 9003 3924
rect 9003 3918 9037 3924
rect 9037 3918 9054 3924
rect 9002 3879 9054 3918
rect 9002 3872 9003 3879
rect 9003 3872 9037 3879
rect 9037 3872 9054 3879
rect 9066 3918 9075 3924
rect 9075 3918 9109 3924
rect 9109 3918 9118 3924
rect 9066 3879 9118 3918
rect 9066 3872 9075 3879
rect 9075 3872 9109 3879
rect 9109 3872 9118 3879
rect 9130 3918 9147 3924
rect 9147 3918 9181 3924
rect 9181 3918 9182 3924
rect 9130 3879 9182 3918
rect 9130 3872 9147 3879
rect 9147 3872 9181 3879
rect 9181 3872 9182 3879
rect 9002 3845 9003 3859
rect 9003 3845 9037 3859
rect 9037 3845 9054 3859
rect 9002 3807 9054 3845
rect 9066 3845 9075 3859
rect 9075 3845 9109 3859
rect 9109 3845 9118 3859
rect 9066 3807 9118 3845
rect 9130 3845 9147 3859
rect 9147 3845 9181 3859
rect 9181 3845 9182 3859
rect 9130 3807 9182 3845
rect 9002 3772 9003 3794
rect 9003 3772 9037 3794
rect 9037 3772 9054 3794
rect 9002 3742 9054 3772
rect 9066 3772 9075 3794
rect 9075 3772 9109 3794
rect 9109 3772 9118 3794
rect 9066 3742 9118 3772
rect 9130 3772 9147 3794
rect 9147 3772 9181 3794
rect 9181 3772 9182 3794
rect 9130 3742 9182 3772
rect 9002 3699 9003 3729
rect 9003 3699 9037 3729
rect 9037 3699 9054 3729
rect 9002 3677 9054 3699
rect 9066 3699 9075 3729
rect 9075 3699 9109 3729
rect 9109 3699 9118 3729
rect 9066 3677 9118 3699
rect 9130 3699 9147 3729
rect 9147 3699 9181 3729
rect 9181 3699 9182 3729
rect 9130 3677 9182 3699
rect 9002 3660 9182 3664
rect 9002 3626 9003 3660
rect 9003 3626 9037 3660
rect 9037 3626 9075 3660
rect 9075 3626 9109 3660
rect 9109 3626 9147 3660
rect 9147 3626 9181 3660
rect 9181 3626 9182 3660
rect 9002 3587 9182 3626
rect 9002 3553 9003 3587
rect 9003 3553 9037 3587
rect 9037 3553 9075 3587
rect 9075 3553 9109 3587
rect 9109 3553 9147 3587
rect 9147 3553 9181 3587
rect 9181 3553 9182 3587
rect 9002 3514 9182 3553
rect 9002 3480 9003 3514
rect 9003 3480 9037 3514
rect 9037 3480 9075 3514
rect 9075 3480 9109 3514
rect 9109 3480 9147 3514
rect 9147 3480 9181 3514
rect 9181 3480 9182 3514
rect 9002 3441 9182 3480
rect 9002 3407 9003 3441
rect 9003 3407 9037 3441
rect 9037 3407 9075 3441
rect 9075 3407 9109 3441
rect 9109 3407 9147 3441
rect 9147 3407 9181 3441
rect 9181 3407 9182 3441
rect 9002 3368 9182 3407
rect 9002 3334 9003 3368
rect 9003 3334 9037 3368
rect 9037 3334 9075 3368
rect 9075 3334 9109 3368
rect 9109 3334 9147 3368
rect 9147 3334 9181 3368
rect 9181 3334 9182 3368
rect 9002 3295 9182 3334
rect 9002 3261 9003 3295
rect 9003 3261 9037 3295
rect 9037 3261 9075 3295
rect 9075 3261 9109 3295
rect 9109 3261 9147 3295
rect 9147 3261 9181 3295
rect 9181 3261 9182 3295
rect 9002 3222 9182 3261
rect 9002 3188 9003 3222
rect 9003 3188 9037 3222
rect 9037 3188 9075 3222
rect 9075 3188 9109 3222
rect 9109 3188 9147 3222
rect 9147 3188 9181 3222
rect 9181 3188 9182 3222
rect 9002 3149 9182 3188
rect 9002 3115 9003 3149
rect 9003 3115 9037 3149
rect 9037 3115 9075 3149
rect 9075 3115 9109 3149
rect 9109 3115 9147 3149
rect 9147 3115 9181 3149
rect 9181 3115 9182 3149
rect 9002 3076 9182 3115
rect 9002 3042 9003 3076
rect 9003 3042 9037 3076
rect 9037 3042 9075 3076
rect 9075 3042 9109 3076
rect 9109 3042 9147 3076
rect 9147 3042 9181 3076
rect 9181 3042 9182 3076
rect 9002 3003 9182 3042
rect 9002 2972 9003 3003
rect 9003 2972 9037 3003
rect 9037 2972 9075 3003
rect 9075 2972 9109 3003
rect 9109 2972 9147 3003
rect 9147 2972 9181 3003
rect 9181 2972 9182 3003
rect 9498 2628 9550 2657
rect 9498 2605 9499 2628
rect 9499 2605 9533 2628
rect 9533 2605 9550 2628
rect 9562 2628 9614 2657
rect 9562 2605 9571 2628
rect 9571 2605 9605 2628
rect 9605 2605 9614 2628
rect 9626 2628 9678 2657
rect 9626 2605 9643 2628
rect 9643 2605 9677 2628
rect 9677 2605 9678 2628
rect 9498 2540 9550 2592
rect 9562 2556 9614 2592
rect 9562 2540 9571 2556
rect 9571 2540 9605 2556
rect 9605 2540 9614 2556
rect 9626 2540 9678 2592
rect 9498 2518 9550 2527
rect 9562 2522 9571 2527
rect 9571 2522 9605 2527
rect 9605 2522 9614 2527
rect 9562 2518 9614 2522
rect 9626 2518 9678 2527
rect 9498 2475 9499 2518
rect 9499 2475 9550 2518
rect 9562 2475 9614 2518
rect 9626 2475 9677 2518
rect 9677 2475 9678 2518
rect 9498 2410 9499 2462
rect 9499 2410 9550 2462
rect 9562 2410 9614 2462
rect 9626 2410 9677 2462
rect 9677 2410 9678 2462
rect 9498 2345 9499 2397
rect 9499 2345 9550 2397
rect 9562 2345 9614 2397
rect 9626 2345 9677 2397
rect 9677 2345 9678 2397
rect 9498 2280 9499 2332
rect 9499 2280 9550 2332
rect 9562 2280 9614 2332
rect 9626 2280 9677 2332
rect 9677 2280 9678 2332
rect 9498 2215 9499 2267
rect 9499 2215 9550 2267
rect 9562 2215 9614 2267
rect 9626 2215 9677 2267
rect 9677 2215 9678 2267
rect 9498 2150 9499 2202
rect 9499 2150 9550 2202
rect 9562 2150 9614 2202
rect 9626 2150 9677 2202
rect 9677 2150 9678 2202
rect 9498 2085 9499 2137
rect 9499 2085 9550 2137
rect 9562 2085 9614 2137
rect 9626 2085 9677 2137
rect 9677 2085 9678 2137
rect 9498 2020 9499 2072
rect 9499 2020 9550 2072
rect 9562 2020 9614 2072
rect 9626 2020 9677 2072
rect 9677 2020 9678 2072
rect 9498 1955 9499 2007
rect 9499 1955 9550 2007
rect 9562 1955 9614 2007
rect 9626 1955 9677 2007
rect 9677 1955 9678 2007
rect 9498 1890 9499 1942
rect 9499 1890 9550 1942
rect 9562 1890 9614 1942
rect 9626 1890 9677 1942
rect 9677 1890 9678 1942
rect 9498 1825 9499 1877
rect 9499 1825 9550 1877
rect 9562 1825 9614 1877
rect 9626 1825 9677 1877
rect 9677 1825 9678 1877
rect 9498 1620 9499 1812
rect 9499 1620 9677 1812
rect 9677 1620 9678 1812
rect 9498 1586 9571 1620
rect 9571 1586 9605 1620
rect 9605 1586 9678 1620
rect 9498 1568 9678 1586
rect 9994 4098 10046 4119
rect 9994 4067 9995 4098
rect 9995 4067 10029 4098
rect 10029 4067 10046 4098
rect 10058 4098 10110 4119
rect 10058 4067 10067 4098
rect 10067 4067 10101 4098
rect 10101 4067 10110 4098
rect 10122 4098 10174 4119
rect 10122 4067 10139 4098
rect 10139 4067 10173 4098
rect 10173 4067 10174 4098
rect 9994 4025 10046 4054
rect 9994 4002 9995 4025
rect 9995 4002 10029 4025
rect 10029 4002 10046 4025
rect 10058 4025 10110 4054
rect 10058 4002 10067 4025
rect 10067 4002 10101 4025
rect 10101 4002 10110 4025
rect 10122 4025 10174 4054
rect 10122 4002 10139 4025
rect 10139 4002 10173 4025
rect 10173 4002 10174 4025
rect 9994 3952 10046 3989
rect 9994 3937 9995 3952
rect 9995 3937 10029 3952
rect 10029 3937 10046 3952
rect 10058 3952 10110 3989
rect 10058 3937 10067 3952
rect 10067 3937 10101 3952
rect 10101 3937 10110 3952
rect 10122 3952 10174 3989
rect 10122 3937 10139 3952
rect 10139 3937 10173 3952
rect 10173 3937 10174 3952
rect 9994 3918 9995 3924
rect 9995 3918 10029 3924
rect 10029 3918 10046 3924
rect 9994 3879 10046 3918
rect 9994 3872 9995 3879
rect 9995 3872 10029 3879
rect 10029 3872 10046 3879
rect 10058 3918 10067 3924
rect 10067 3918 10101 3924
rect 10101 3918 10110 3924
rect 10058 3879 10110 3918
rect 10058 3872 10067 3879
rect 10067 3872 10101 3879
rect 10101 3872 10110 3879
rect 10122 3918 10139 3924
rect 10139 3918 10173 3924
rect 10173 3918 10174 3924
rect 10122 3879 10174 3918
rect 10122 3872 10139 3879
rect 10139 3872 10173 3879
rect 10173 3872 10174 3879
rect 9994 3845 9995 3859
rect 9995 3845 10029 3859
rect 10029 3845 10046 3859
rect 9994 3807 10046 3845
rect 10058 3845 10067 3859
rect 10067 3845 10101 3859
rect 10101 3845 10110 3859
rect 10058 3807 10110 3845
rect 10122 3845 10139 3859
rect 10139 3845 10173 3859
rect 10173 3845 10174 3859
rect 10122 3807 10174 3845
rect 9994 3772 9995 3794
rect 9995 3772 10029 3794
rect 10029 3772 10046 3794
rect 9994 3742 10046 3772
rect 10058 3772 10067 3794
rect 10067 3772 10101 3794
rect 10101 3772 10110 3794
rect 10058 3742 10110 3772
rect 10122 3772 10139 3794
rect 10139 3772 10173 3794
rect 10173 3772 10174 3794
rect 10122 3742 10174 3772
rect 9994 3699 9995 3729
rect 9995 3699 10029 3729
rect 10029 3699 10046 3729
rect 9994 3677 10046 3699
rect 10058 3699 10067 3729
rect 10067 3699 10101 3729
rect 10101 3699 10110 3729
rect 10058 3677 10110 3699
rect 10122 3699 10139 3729
rect 10139 3699 10173 3729
rect 10173 3699 10174 3729
rect 10122 3677 10174 3699
rect 9994 3660 10174 3664
rect 9994 3626 9995 3660
rect 9995 3626 10029 3660
rect 10029 3626 10067 3660
rect 10067 3626 10101 3660
rect 10101 3626 10139 3660
rect 10139 3626 10173 3660
rect 10173 3626 10174 3660
rect 9994 3587 10174 3626
rect 9994 3553 9995 3587
rect 9995 3553 10029 3587
rect 10029 3553 10067 3587
rect 10067 3553 10101 3587
rect 10101 3553 10139 3587
rect 10139 3553 10173 3587
rect 10173 3553 10174 3587
rect 9994 3514 10174 3553
rect 9994 3480 9995 3514
rect 9995 3480 10029 3514
rect 10029 3480 10067 3514
rect 10067 3480 10101 3514
rect 10101 3480 10139 3514
rect 10139 3480 10173 3514
rect 10173 3480 10174 3514
rect 9994 3441 10174 3480
rect 9994 3407 9995 3441
rect 9995 3407 10029 3441
rect 10029 3407 10067 3441
rect 10067 3407 10101 3441
rect 10101 3407 10139 3441
rect 10139 3407 10173 3441
rect 10173 3407 10174 3441
rect 9994 3368 10174 3407
rect 9994 3334 9995 3368
rect 9995 3334 10029 3368
rect 10029 3334 10067 3368
rect 10067 3334 10101 3368
rect 10101 3334 10139 3368
rect 10139 3334 10173 3368
rect 10173 3334 10174 3368
rect 9994 3295 10174 3334
rect 9994 3261 9995 3295
rect 9995 3261 10029 3295
rect 10029 3261 10067 3295
rect 10067 3261 10101 3295
rect 10101 3261 10139 3295
rect 10139 3261 10173 3295
rect 10173 3261 10174 3295
rect 9994 3222 10174 3261
rect 9994 3188 9995 3222
rect 9995 3188 10029 3222
rect 10029 3188 10067 3222
rect 10067 3188 10101 3222
rect 10101 3188 10139 3222
rect 10139 3188 10173 3222
rect 10173 3188 10174 3222
rect 9994 3149 10174 3188
rect 9994 3115 9995 3149
rect 9995 3115 10029 3149
rect 10029 3115 10067 3149
rect 10067 3115 10101 3149
rect 10101 3115 10139 3149
rect 10139 3115 10173 3149
rect 10173 3115 10174 3149
rect 9994 3076 10174 3115
rect 9994 3042 9995 3076
rect 9995 3042 10029 3076
rect 10029 3042 10067 3076
rect 10067 3042 10101 3076
rect 10101 3042 10139 3076
rect 10139 3042 10173 3076
rect 10173 3042 10174 3076
rect 9994 3003 10174 3042
rect 9994 2972 9995 3003
rect 9995 2972 10029 3003
rect 10029 2972 10067 3003
rect 10067 2972 10101 3003
rect 10101 2972 10139 3003
rect 10139 2972 10173 3003
rect 10173 2972 10174 3003
rect 10490 2628 10542 2657
rect 10490 2605 10491 2628
rect 10491 2605 10525 2628
rect 10525 2605 10542 2628
rect 10554 2628 10606 2657
rect 10554 2605 10563 2628
rect 10563 2605 10597 2628
rect 10597 2605 10606 2628
rect 10618 2628 10670 2657
rect 10618 2605 10635 2628
rect 10635 2605 10669 2628
rect 10669 2605 10670 2628
rect 10490 2540 10542 2592
rect 10554 2556 10606 2592
rect 10554 2540 10563 2556
rect 10563 2540 10597 2556
rect 10597 2540 10606 2556
rect 10618 2540 10670 2592
rect 10490 2518 10542 2527
rect 10554 2522 10563 2527
rect 10563 2522 10597 2527
rect 10597 2522 10606 2527
rect 10554 2518 10606 2522
rect 10618 2518 10670 2527
rect 10490 2475 10491 2518
rect 10491 2475 10542 2518
rect 10554 2475 10606 2518
rect 10618 2475 10669 2518
rect 10669 2475 10670 2518
rect 10490 2410 10491 2462
rect 10491 2410 10542 2462
rect 10554 2410 10606 2462
rect 10618 2410 10669 2462
rect 10669 2410 10670 2462
rect 10490 2345 10491 2397
rect 10491 2345 10542 2397
rect 10554 2345 10606 2397
rect 10618 2345 10669 2397
rect 10669 2345 10670 2397
rect 10490 2280 10491 2332
rect 10491 2280 10542 2332
rect 10554 2280 10606 2332
rect 10618 2280 10669 2332
rect 10669 2280 10670 2332
rect 10490 2215 10491 2267
rect 10491 2215 10542 2267
rect 10554 2215 10606 2267
rect 10618 2215 10669 2267
rect 10669 2215 10670 2267
rect 10490 2150 10491 2202
rect 10491 2150 10542 2202
rect 10554 2150 10606 2202
rect 10618 2150 10669 2202
rect 10669 2150 10670 2202
rect 10490 2085 10491 2137
rect 10491 2085 10542 2137
rect 10554 2085 10606 2137
rect 10618 2085 10669 2137
rect 10669 2085 10670 2137
rect 10490 2020 10491 2072
rect 10491 2020 10542 2072
rect 10554 2020 10606 2072
rect 10618 2020 10669 2072
rect 10669 2020 10670 2072
rect 10490 1955 10491 2007
rect 10491 1955 10542 2007
rect 10554 1955 10606 2007
rect 10618 1955 10669 2007
rect 10669 1955 10670 2007
rect 10490 1890 10491 1942
rect 10491 1890 10542 1942
rect 10554 1890 10606 1942
rect 10618 1890 10669 1942
rect 10669 1890 10670 1942
rect 10490 1825 10491 1877
rect 10491 1825 10542 1877
rect 10554 1825 10606 1877
rect 10618 1825 10669 1877
rect 10669 1825 10670 1877
rect 10490 1620 10491 1812
rect 10491 1620 10669 1812
rect 10669 1620 10670 1812
rect 10490 1586 10563 1620
rect 10563 1586 10597 1620
rect 10597 1586 10670 1620
rect 10490 1568 10670 1586
rect 10986 4098 11038 4119
rect 10986 4067 10987 4098
rect 10987 4067 11021 4098
rect 11021 4067 11038 4098
rect 11050 4098 11102 4119
rect 11050 4067 11059 4098
rect 11059 4067 11093 4098
rect 11093 4067 11102 4098
rect 11114 4098 11166 4119
rect 11114 4067 11131 4098
rect 11131 4067 11165 4098
rect 11165 4067 11166 4098
rect 10986 4025 11038 4054
rect 10986 4002 10987 4025
rect 10987 4002 11021 4025
rect 11021 4002 11038 4025
rect 11050 4025 11102 4054
rect 11050 4002 11059 4025
rect 11059 4002 11093 4025
rect 11093 4002 11102 4025
rect 11114 4025 11166 4054
rect 11114 4002 11131 4025
rect 11131 4002 11165 4025
rect 11165 4002 11166 4025
rect 10986 3952 11038 3989
rect 10986 3937 10987 3952
rect 10987 3937 11021 3952
rect 11021 3937 11038 3952
rect 11050 3952 11102 3989
rect 11050 3937 11059 3952
rect 11059 3937 11093 3952
rect 11093 3937 11102 3952
rect 11114 3952 11166 3989
rect 11114 3937 11131 3952
rect 11131 3937 11165 3952
rect 11165 3937 11166 3952
rect 10986 3918 10987 3924
rect 10987 3918 11021 3924
rect 11021 3918 11038 3924
rect 10986 3879 11038 3918
rect 10986 3872 10987 3879
rect 10987 3872 11021 3879
rect 11021 3872 11038 3879
rect 11050 3918 11059 3924
rect 11059 3918 11093 3924
rect 11093 3918 11102 3924
rect 11050 3879 11102 3918
rect 11050 3872 11059 3879
rect 11059 3872 11093 3879
rect 11093 3872 11102 3879
rect 11114 3918 11131 3924
rect 11131 3918 11165 3924
rect 11165 3918 11166 3924
rect 11114 3879 11166 3918
rect 11114 3872 11131 3879
rect 11131 3872 11165 3879
rect 11165 3872 11166 3879
rect 10986 3845 10987 3859
rect 10987 3845 11021 3859
rect 11021 3845 11038 3859
rect 10986 3807 11038 3845
rect 11050 3845 11059 3859
rect 11059 3845 11093 3859
rect 11093 3845 11102 3859
rect 11050 3807 11102 3845
rect 11114 3845 11131 3859
rect 11131 3845 11165 3859
rect 11165 3845 11166 3859
rect 11114 3807 11166 3845
rect 10986 3772 10987 3794
rect 10987 3772 11021 3794
rect 11021 3772 11038 3794
rect 10986 3742 11038 3772
rect 11050 3772 11059 3794
rect 11059 3772 11093 3794
rect 11093 3772 11102 3794
rect 11050 3742 11102 3772
rect 11114 3772 11131 3794
rect 11131 3772 11165 3794
rect 11165 3772 11166 3794
rect 11114 3742 11166 3772
rect 10986 3699 10987 3729
rect 10987 3699 11021 3729
rect 11021 3699 11038 3729
rect 10986 3677 11038 3699
rect 11050 3699 11059 3729
rect 11059 3699 11093 3729
rect 11093 3699 11102 3729
rect 11050 3677 11102 3699
rect 11114 3699 11131 3729
rect 11131 3699 11165 3729
rect 11165 3699 11166 3729
rect 11114 3677 11166 3699
rect 10986 3660 11166 3664
rect 10986 3626 10987 3660
rect 10987 3626 11021 3660
rect 11021 3626 11059 3660
rect 11059 3626 11093 3660
rect 11093 3626 11131 3660
rect 11131 3626 11165 3660
rect 11165 3626 11166 3660
rect 10986 3587 11166 3626
rect 10986 3553 10987 3587
rect 10987 3553 11021 3587
rect 11021 3553 11059 3587
rect 11059 3553 11093 3587
rect 11093 3553 11131 3587
rect 11131 3553 11165 3587
rect 11165 3553 11166 3587
rect 10986 3514 11166 3553
rect 10986 3480 10987 3514
rect 10987 3480 11021 3514
rect 11021 3480 11059 3514
rect 11059 3480 11093 3514
rect 11093 3480 11131 3514
rect 11131 3480 11165 3514
rect 11165 3480 11166 3514
rect 10986 3441 11166 3480
rect 10986 3407 10987 3441
rect 10987 3407 11021 3441
rect 11021 3407 11059 3441
rect 11059 3407 11093 3441
rect 11093 3407 11131 3441
rect 11131 3407 11165 3441
rect 11165 3407 11166 3441
rect 10986 3368 11166 3407
rect 10986 3334 10987 3368
rect 10987 3334 11021 3368
rect 11021 3334 11059 3368
rect 11059 3334 11093 3368
rect 11093 3334 11131 3368
rect 11131 3334 11165 3368
rect 11165 3334 11166 3368
rect 10986 3295 11166 3334
rect 10986 3261 10987 3295
rect 10987 3261 11021 3295
rect 11021 3261 11059 3295
rect 11059 3261 11093 3295
rect 11093 3261 11131 3295
rect 11131 3261 11165 3295
rect 11165 3261 11166 3295
rect 10986 3222 11166 3261
rect 10986 3188 10987 3222
rect 10987 3188 11021 3222
rect 11021 3188 11059 3222
rect 11059 3188 11093 3222
rect 11093 3188 11131 3222
rect 11131 3188 11165 3222
rect 11165 3188 11166 3222
rect 10986 3149 11166 3188
rect 10986 3115 10987 3149
rect 10987 3115 11021 3149
rect 11021 3115 11059 3149
rect 11059 3115 11093 3149
rect 11093 3115 11131 3149
rect 11131 3115 11165 3149
rect 11165 3115 11166 3149
rect 10986 3076 11166 3115
rect 10986 3042 10987 3076
rect 10987 3042 11021 3076
rect 11021 3042 11059 3076
rect 11059 3042 11093 3076
rect 11093 3042 11131 3076
rect 11131 3042 11165 3076
rect 11165 3042 11166 3076
rect 10986 3003 11166 3042
rect 10986 2972 10987 3003
rect 10987 2972 11021 3003
rect 11021 2972 11059 3003
rect 11059 2972 11093 3003
rect 11093 2972 11131 3003
rect 11131 2972 11165 3003
rect 11165 2972 11166 3003
rect 11482 2628 11534 2657
rect 11482 2605 11483 2628
rect 11483 2605 11517 2628
rect 11517 2605 11534 2628
rect 11546 2628 11598 2657
rect 11546 2605 11555 2628
rect 11555 2605 11589 2628
rect 11589 2605 11598 2628
rect 11610 2628 11662 2657
rect 11610 2605 11627 2628
rect 11627 2605 11661 2628
rect 11661 2605 11662 2628
rect 11482 2540 11534 2592
rect 11546 2556 11598 2592
rect 11546 2540 11555 2556
rect 11555 2540 11589 2556
rect 11589 2540 11598 2556
rect 11610 2540 11662 2592
rect 11482 2518 11534 2527
rect 11546 2522 11555 2527
rect 11555 2522 11589 2527
rect 11589 2522 11598 2527
rect 11546 2518 11598 2522
rect 11610 2518 11662 2527
rect 11482 2475 11483 2518
rect 11483 2475 11534 2518
rect 11546 2475 11598 2518
rect 11610 2475 11661 2518
rect 11661 2475 11662 2518
rect 11482 2410 11483 2462
rect 11483 2410 11534 2462
rect 11546 2410 11598 2462
rect 11610 2410 11661 2462
rect 11661 2410 11662 2462
rect 11482 2345 11483 2397
rect 11483 2345 11534 2397
rect 11546 2345 11598 2397
rect 11610 2345 11661 2397
rect 11661 2345 11662 2397
rect 11482 2280 11483 2332
rect 11483 2280 11534 2332
rect 11546 2280 11598 2332
rect 11610 2280 11661 2332
rect 11661 2280 11662 2332
rect 11482 2215 11483 2267
rect 11483 2215 11534 2267
rect 11546 2215 11598 2267
rect 11610 2215 11661 2267
rect 11661 2215 11662 2267
rect 11482 2150 11483 2202
rect 11483 2150 11534 2202
rect 11546 2150 11598 2202
rect 11610 2150 11661 2202
rect 11661 2150 11662 2202
rect 11482 2085 11483 2137
rect 11483 2085 11534 2137
rect 11546 2085 11598 2137
rect 11610 2085 11661 2137
rect 11661 2085 11662 2137
rect 11482 2020 11483 2072
rect 11483 2020 11534 2072
rect 11546 2020 11598 2072
rect 11610 2020 11661 2072
rect 11661 2020 11662 2072
rect 11482 1955 11483 2007
rect 11483 1955 11534 2007
rect 11546 1955 11598 2007
rect 11610 1955 11661 2007
rect 11661 1955 11662 2007
rect 11482 1890 11483 1942
rect 11483 1890 11534 1942
rect 11546 1890 11598 1942
rect 11610 1890 11661 1942
rect 11661 1890 11662 1942
rect 11482 1825 11483 1877
rect 11483 1825 11534 1877
rect 11546 1825 11598 1877
rect 11610 1825 11661 1877
rect 11661 1825 11662 1877
rect 11482 1620 11483 1812
rect 11483 1620 11661 1812
rect 11661 1620 11662 1812
rect 11482 1586 11555 1620
rect 11555 1586 11589 1620
rect 11589 1586 11662 1620
rect 11482 1568 11662 1586
rect 11978 4098 12030 4119
rect 11978 4067 11979 4098
rect 11979 4067 12013 4098
rect 12013 4067 12030 4098
rect 12042 4098 12094 4119
rect 12042 4067 12051 4098
rect 12051 4067 12085 4098
rect 12085 4067 12094 4098
rect 12106 4098 12158 4119
rect 12106 4067 12123 4098
rect 12123 4067 12157 4098
rect 12157 4067 12158 4098
rect 11978 4025 12030 4054
rect 11978 4002 11979 4025
rect 11979 4002 12013 4025
rect 12013 4002 12030 4025
rect 12042 4025 12094 4054
rect 12042 4002 12051 4025
rect 12051 4002 12085 4025
rect 12085 4002 12094 4025
rect 12106 4025 12158 4054
rect 12106 4002 12123 4025
rect 12123 4002 12157 4025
rect 12157 4002 12158 4025
rect 11978 3952 12030 3989
rect 11978 3937 11979 3952
rect 11979 3937 12013 3952
rect 12013 3937 12030 3952
rect 12042 3952 12094 3989
rect 12042 3937 12051 3952
rect 12051 3937 12085 3952
rect 12085 3937 12094 3952
rect 12106 3952 12158 3989
rect 12106 3937 12123 3952
rect 12123 3937 12157 3952
rect 12157 3937 12158 3952
rect 11978 3918 11979 3924
rect 11979 3918 12013 3924
rect 12013 3918 12030 3924
rect 11978 3879 12030 3918
rect 11978 3872 11979 3879
rect 11979 3872 12013 3879
rect 12013 3872 12030 3879
rect 12042 3918 12051 3924
rect 12051 3918 12085 3924
rect 12085 3918 12094 3924
rect 12042 3879 12094 3918
rect 12042 3872 12051 3879
rect 12051 3872 12085 3879
rect 12085 3872 12094 3879
rect 12106 3918 12123 3924
rect 12123 3918 12157 3924
rect 12157 3918 12158 3924
rect 12106 3879 12158 3918
rect 12106 3872 12123 3879
rect 12123 3872 12157 3879
rect 12157 3872 12158 3879
rect 11978 3845 11979 3859
rect 11979 3845 12013 3859
rect 12013 3845 12030 3859
rect 11978 3807 12030 3845
rect 12042 3845 12051 3859
rect 12051 3845 12085 3859
rect 12085 3845 12094 3859
rect 12042 3807 12094 3845
rect 12106 3845 12123 3859
rect 12123 3845 12157 3859
rect 12157 3845 12158 3859
rect 12106 3807 12158 3845
rect 11978 3772 11979 3794
rect 11979 3772 12013 3794
rect 12013 3772 12030 3794
rect 11978 3742 12030 3772
rect 12042 3772 12051 3794
rect 12051 3772 12085 3794
rect 12085 3772 12094 3794
rect 12042 3742 12094 3772
rect 12106 3772 12123 3794
rect 12123 3772 12157 3794
rect 12157 3772 12158 3794
rect 12106 3742 12158 3772
rect 11978 3699 11979 3729
rect 11979 3699 12013 3729
rect 12013 3699 12030 3729
rect 11978 3677 12030 3699
rect 12042 3699 12051 3729
rect 12051 3699 12085 3729
rect 12085 3699 12094 3729
rect 12042 3677 12094 3699
rect 12106 3699 12123 3729
rect 12123 3699 12157 3729
rect 12157 3699 12158 3729
rect 12106 3677 12158 3699
rect 11978 3660 12158 3664
rect 11978 3626 11979 3660
rect 11979 3626 12013 3660
rect 12013 3626 12051 3660
rect 12051 3626 12085 3660
rect 12085 3626 12123 3660
rect 12123 3626 12157 3660
rect 12157 3626 12158 3660
rect 11978 3587 12158 3626
rect 11978 3553 11979 3587
rect 11979 3553 12013 3587
rect 12013 3553 12051 3587
rect 12051 3553 12085 3587
rect 12085 3553 12123 3587
rect 12123 3553 12157 3587
rect 12157 3553 12158 3587
rect 11978 3514 12158 3553
rect 11978 3480 11979 3514
rect 11979 3480 12013 3514
rect 12013 3480 12051 3514
rect 12051 3480 12085 3514
rect 12085 3480 12123 3514
rect 12123 3480 12157 3514
rect 12157 3480 12158 3514
rect 11978 3441 12158 3480
rect 11978 3407 11979 3441
rect 11979 3407 12013 3441
rect 12013 3407 12051 3441
rect 12051 3407 12085 3441
rect 12085 3407 12123 3441
rect 12123 3407 12157 3441
rect 12157 3407 12158 3441
rect 11978 3368 12158 3407
rect 11978 3334 11979 3368
rect 11979 3334 12013 3368
rect 12013 3334 12051 3368
rect 12051 3334 12085 3368
rect 12085 3334 12123 3368
rect 12123 3334 12157 3368
rect 12157 3334 12158 3368
rect 11978 3295 12158 3334
rect 11978 3261 11979 3295
rect 11979 3261 12013 3295
rect 12013 3261 12051 3295
rect 12051 3261 12085 3295
rect 12085 3261 12123 3295
rect 12123 3261 12157 3295
rect 12157 3261 12158 3295
rect 11978 3222 12158 3261
rect 11978 3188 11979 3222
rect 11979 3188 12013 3222
rect 12013 3188 12051 3222
rect 12051 3188 12085 3222
rect 12085 3188 12123 3222
rect 12123 3188 12157 3222
rect 12157 3188 12158 3222
rect 11978 3149 12158 3188
rect 11978 3115 11979 3149
rect 11979 3115 12013 3149
rect 12013 3115 12051 3149
rect 12051 3115 12085 3149
rect 12085 3115 12123 3149
rect 12123 3115 12157 3149
rect 12157 3115 12158 3149
rect 11978 3076 12158 3115
rect 11978 3042 11979 3076
rect 11979 3042 12013 3076
rect 12013 3042 12051 3076
rect 12051 3042 12085 3076
rect 12085 3042 12123 3076
rect 12123 3042 12157 3076
rect 12157 3042 12158 3076
rect 11978 3003 12158 3042
rect 11978 2972 11979 3003
rect 11979 2972 12013 3003
rect 12013 2972 12051 3003
rect 12051 2972 12085 3003
rect 12085 2972 12123 3003
rect 12123 2972 12157 3003
rect 12157 2972 12158 3003
rect 12474 2628 12526 2657
rect 12474 2605 12475 2628
rect 12475 2605 12509 2628
rect 12509 2605 12526 2628
rect 12538 2628 12590 2657
rect 12538 2605 12547 2628
rect 12547 2605 12581 2628
rect 12581 2605 12590 2628
rect 12602 2628 12654 2657
rect 12602 2605 12619 2628
rect 12619 2605 12653 2628
rect 12653 2605 12654 2628
rect 12474 2540 12526 2592
rect 12538 2556 12590 2592
rect 12538 2540 12547 2556
rect 12547 2540 12581 2556
rect 12581 2540 12590 2556
rect 12602 2540 12654 2592
rect 12474 2518 12526 2527
rect 12538 2522 12547 2527
rect 12547 2522 12581 2527
rect 12581 2522 12590 2527
rect 12538 2518 12590 2522
rect 12602 2518 12654 2527
rect 12474 2475 12475 2518
rect 12475 2475 12526 2518
rect 12538 2475 12590 2518
rect 12602 2475 12653 2518
rect 12653 2475 12654 2518
rect 12474 2410 12475 2462
rect 12475 2410 12526 2462
rect 12538 2410 12590 2462
rect 12602 2410 12653 2462
rect 12653 2410 12654 2462
rect 12474 2345 12475 2397
rect 12475 2345 12526 2397
rect 12538 2345 12590 2397
rect 12602 2345 12653 2397
rect 12653 2345 12654 2397
rect 12474 2280 12475 2332
rect 12475 2280 12526 2332
rect 12538 2280 12590 2332
rect 12602 2280 12653 2332
rect 12653 2280 12654 2332
rect 12474 2215 12475 2267
rect 12475 2215 12526 2267
rect 12538 2215 12590 2267
rect 12602 2215 12653 2267
rect 12653 2215 12654 2267
rect 12474 2150 12475 2202
rect 12475 2150 12526 2202
rect 12538 2150 12590 2202
rect 12602 2150 12653 2202
rect 12653 2150 12654 2202
rect 12474 2085 12475 2137
rect 12475 2085 12526 2137
rect 12538 2085 12590 2137
rect 12602 2085 12653 2137
rect 12653 2085 12654 2137
rect 12474 2020 12475 2072
rect 12475 2020 12526 2072
rect 12538 2020 12590 2072
rect 12602 2020 12653 2072
rect 12653 2020 12654 2072
rect 12474 1955 12475 2007
rect 12475 1955 12526 2007
rect 12538 1955 12590 2007
rect 12602 1955 12653 2007
rect 12653 1955 12654 2007
rect 12474 1890 12475 1942
rect 12475 1890 12526 1942
rect 12538 1890 12590 1942
rect 12602 1890 12653 1942
rect 12653 1890 12654 1942
rect 12474 1825 12475 1877
rect 12475 1825 12526 1877
rect 12538 1825 12590 1877
rect 12602 1825 12653 1877
rect 12653 1825 12654 1877
rect 12474 1620 12475 1812
rect 12475 1620 12653 1812
rect 12653 1620 12654 1812
rect 12474 1586 12547 1620
rect 12547 1586 12581 1620
rect 12581 1586 12654 1620
rect 12474 1568 12654 1586
rect 12970 4098 13022 4119
rect 12970 4067 12971 4098
rect 12971 4067 13005 4098
rect 13005 4067 13022 4098
rect 13034 4098 13086 4119
rect 13034 4067 13043 4098
rect 13043 4067 13077 4098
rect 13077 4067 13086 4098
rect 13098 4098 13150 4119
rect 13098 4067 13115 4098
rect 13115 4067 13149 4098
rect 13149 4067 13150 4098
rect 12970 4025 13022 4054
rect 12970 4002 12971 4025
rect 12971 4002 13005 4025
rect 13005 4002 13022 4025
rect 13034 4025 13086 4054
rect 13034 4002 13043 4025
rect 13043 4002 13077 4025
rect 13077 4002 13086 4025
rect 13098 4025 13150 4054
rect 13098 4002 13115 4025
rect 13115 4002 13149 4025
rect 13149 4002 13150 4025
rect 12970 3952 13022 3989
rect 12970 3937 12971 3952
rect 12971 3937 13005 3952
rect 13005 3937 13022 3952
rect 13034 3952 13086 3989
rect 13034 3937 13043 3952
rect 13043 3937 13077 3952
rect 13077 3937 13086 3952
rect 13098 3952 13150 3989
rect 13098 3937 13115 3952
rect 13115 3937 13149 3952
rect 13149 3937 13150 3952
rect 12970 3918 12971 3924
rect 12971 3918 13005 3924
rect 13005 3918 13022 3924
rect 12970 3879 13022 3918
rect 12970 3872 12971 3879
rect 12971 3872 13005 3879
rect 13005 3872 13022 3879
rect 13034 3918 13043 3924
rect 13043 3918 13077 3924
rect 13077 3918 13086 3924
rect 13034 3879 13086 3918
rect 13034 3872 13043 3879
rect 13043 3872 13077 3879
rect 13077 3872 13086 3879
rect 13098 3918 13115 3924
rect 13115 3918 13149 3924
rect 13149 3918 13150 3924
rect 13098 3879 13150 3918
rect 13098 3872 13115 3879
rect 13115 3872 13149 3879
rect 13149 3872 13150 3879
rect 12970 3845 12971 3859
rect 12971 3845 13005 3859
rect 13005 3845 13022 3859
rect 12970 3807 13022 3845
rect 13034 3845 13043 3859
rect 13043 3845 13077 3859
rect 13077 3845 13086 3859
rect 13034 3807 13086 3845
rect 13098 3845 13115 3859
rect 13115 3845 13149 3859
rect 13149 3845 13150 3859
rect 13098 3807 13150 3845
rect 12970 3772 12971 3794
rect 12971 3772 13005 3794
rect 13005 3772 13022 3794
rect 12970 3742 13022 3772
rect 13034 3772 13043 3794
rect 13043 3772 13077 3794
rect 13077 3772 13086 3794
rect 13034 3742 13086 3772
rect 13098 3772 13115 3794
rect 13115 3772 13149 3794
rect 13149 3772 13150 3794
rect 13098 3742 13150 3772
rect 12970 3699 12971 3729
rect 12971 3699 13005 3729
rect 13005 3699 13022 3729
rect 12970 3677 13022 3699
rect 13034 3699 13043 3729
rect 13043 3699 13077 3729
rect 13077 3699 13086 3729
rect 13034 3677 13086 3699
rect 13098 3699 13115 3729
rect 13115 3699 13149 3729
rect 13149 3699 13150 3729
rect 13098 3677 13150 3699
rect 12970 3660 13150 3664
rect 12970 3626 12971 3660
rect 12971 3626 13005 3660
rect 13005 3626 13043 3660
rect 13043 3626 13077 3660
rect 13077 3626 13115 3660
rect 13115 3626 13149 3660
rect 13149 3626 13150 3660
rect 12970 3587 13150 3626
rect 12970 3553 12971 3587
rect 12971 3553 13005 3587
rect 13005 3553 13043 3587
rect 13043 3553 13077 3587
rect 13077 3553 13115 3587
rect 13115 3553 13149 3587
rect 13149 3553 13150 3587
rect 12970 3514 13150 3553
rect 12970 3480 12971 3514
rect 12971 3480 13005 3514
rect 13005 3480 13043 3514
rect 13043 3480 13077 3514
rect 13077 3480 13115 3514
rect 13115 3480 13149 3514
rect 13149 3480 13150 3514
rect 12970 3441 13150 3480
rect 12970 3407 12971 3441
rect 12971 3407 13005 3441
rect 13005 3407 13043 3441
rect 13043 3407 13077 3441
rect 13077 3407 13115 3441
rect 13115 3407 13149 3441
rect 13149 3407 13150 3441
rect 12970 3368 13150 3407
rect 12970 3334 12971 3368
rect 12971 3334 13005 3368
rect 13005 3334 13043 3368
rect 13043 3334 13077 3368
rect 13077 3334 13115 3368
rect 13115 3334 13149 3368
rect 13149 3334 13150 3368
rect 12970 3295 13150 3334
rect 12970 3261 12971 3295
rect 12971 3261 13005 3295
rect 13005 3261 13043 3295
rect 13043 3261 13077 3295
rect 13077 3261 13115 3295
rect 13115 3261 13149 3295
rect 13149 3261 13150 3295
rect 12970 3222 13150 3261
rect 12970 3188 12971 3222
rect 12971 3188 13005 3222
rect 13005 3188 13043 3222
rect 13043 3188 13077 3222
rect 13077 3188 13115 3222
rect 13115 3188 13149 3222
rect 13149 3188 13150 3222
rect 12970 3149 13150 3188
rect 12970 3115 12971 3149
rect 12971 3115 13005 3149
rect 13005 3115 13043 3149
rect 13043 3115 13077 3149
rect 13077 3115 13115 3149
rect 13115 3115 13149 3149
rect 13149 3115 13150 3149
rect 12970 3076 13150 3115
rect 12970 3042 12971 3076
rect 12971 3042 13005 3076
rect 13005 3042 13043 3076
rect 13043 3042 13077 3076
rect 13077 3042 13115 3076
rect 13115 3042 13149 3076
rect 13149 3042 13150 3076
rect 12970 3003 13150 3042
rect 12970 2972 12971 3003
rect 12971 2972 13005 3003
rect 13005 2972 13043 3003
rect 13043 2972 13077 3003
rect 13077 2972 13115 3003
rect 13115 2972 13149 3003
rect 13149 2972 13150 3003
rect 13466 2628 13518 2657
rect 13466 2605 13467 2628
rect 13467 2605 13501 2628
rect 13501 2605 13518 2628
rect 13530 2628 13582 2657
rect 13530 2605 13539 2628
rect 13539 2605 13573 2628
rect 13573 2605 13582 2628
rect 13594 2628 13646 2657
rect 13594 2605 13611 2628
rect 13611 2605 13645 2628
rect 13645 2605 13646 2628
rect 13466 2540 13518 2592
rect 13530 2556 13582 2592
rect 13530 2540 13539 2556
rect 13539 2540 13573 2556
rect 13573 2540 13582 2556
rect 13594 2540 13646 2592
rect 13466 2518 13518 2527
rect 13530 2522 13539 2527
rect 13539 2522 13573 2527
rect 13573 2522 13582 2527
rect 13530 2518 13582 2522
rect 13594 2518 13646 2527
rect 13466 2475 13467 2518
rect 13467 2475 13518 2518
rect 13530 2475 13582 2518
rect 13594 2475 13645 2518
rect 13645 2475 13646 2518
rect 13466 2410 13467 2462
rect 13467 2410 13518 2462
rect 13530 2410 13582 2462
rect 13594 2410 13645 2462
rect 13645 2410 13646 2462
rect 13466 2345 13467 2397
rect 13467 2345 13518 2397
rect 13530 2345 13582 2397
rect 13594 2345 13645 2397
rect 13645 2345 13646 2397
rect 13466 2280 13467 2332
rect 13467 2280 13518 2332
rect 13530 2280 13582 2332
rect 13594 2280 13645 2332
rect 13645 2280 13646 2332
rect 13466 2215 13467 2267
rect 13467 2215 13518 2267
rect 13530 2215 13582 2267
rect 13594 2215 13645 2267
rect 13645 2215 13646 2267
rect 13466 2150 13467 2202
rect 13467 2150 13518 2202
rect 13530 2150 13582 2202
rect 13594 2150 13645 2202
rect 13645 2150 13646 2202
rect 13466 2085 13467 2137
rect 13467 2085 13518 2137
rect 13530 2085 13582 2137
rect 13594 2085 13645 2137
rect 13645 2085 13646 2137
rect 13466 2020 13467 2072
rect 13467 2020 13518 2072
rect 13530 2020 13582 2072
rect 13594 2020 13645 2072
rect 13645 2020 13646 2072
rect 13466 1955 13467 2007
rect 13467 1955 13518 2007
rect 13530 1955 13582 2007
rect 13594 1955 13645 2007
rect 13645 1955 13646 2007
rect 13466 1890 13467 1942
rect 13467 1890 13518 1942
rect 13530 1890 13582 1942
rect 13594 1890 13645 1942
rect 13645 1890 13646 1942
rect 13466 1825 13467 1877
rect 13467 1825 13518 1877
rect 13530 1825 13582 1877
rect 13594 1825 13645 1877
rect 13645 1825 13646 1877
rect 13466 1620 13467 1812
rect 13467 1620 13645 1812
rect 13645 1620 13646 1812
rect 13466 1586 13539 1620
rect 13539 1586 13573 1620
rect 13573 1586 13646 1620
rect 13466 1568 13646 1586
rect 13990 4098 14042 4119
rect 13990 4067 13999 4098
rect 13999 4067 14033 4098
rect 14033 4067 14042 4098
rect 14062 4067 14114 4119
rect 13990 4025 14042 4055
rect 13990 4003 13999 4025
rect 13999 4003 14033 4025
rect 14033 4003 14042 4025
rect 14062 4003 14114 4055
rect 13990 3952 14042 3991
rect 13990 3939 13999 3952
rect 13999 3939 14033 3952
rect 14033 3939 14042 3952
rect 14062 3939 14114 3991
rect 13990 3918 13999 3927
rect 13999 3918 14033 3927
rect 14033 3918 14042 3927
rect 13990 3879 14042 3918
rect 13990 3875 13999 3879
rect 13999 3875 14033 3879
rect 14033 3875 14042 3879
rect 14062 3875 14114 3927
rect 13990 3845 13999 3863
rect 13999 3845 14033 3863
rect 14033 3845 14042 3863
rect 13990 3811 14042 3845
rect 14062 3811 14114 3863
rect 13990 3772 13999 3799
rect 13999 3772 14033 3799
rect 14033 3772 14042 3799
rect 13990 3747 14042 3772
rect 14062 3747 14114 3799
rect 13990 3733 14042 3735
rect 13990 3699 13999 3733
rect 13999 3699 14033 3733
rect 14033 3699 14042 3733
rect 13990 3683 14042 3699
rect 14062 3683 14114 3735
rect 13990 3660 14042 3671
rect 13990 3626 13999 3660
rect 13999 3626 14033 3660
rect 14033 3626 14042 3660
rect 13990 3619 14042 3626
rect 14062 3619 14114 3671
rect 13990 3587 14042 3607
rect 13990 3555 13999 3587
rect 13999 3555 14033 3587
rect 14033 3555 14042 3587
rect 14062 3555 14114 3607
rect 13990 3514 14042 3543
rect 13990 3491 13999 3514
rect 13999 3491 14033 3514
rect 14033 3491 14042 3514
rect 14062 3491 14114 3543
rect 13990 3441 14042 3479
rect 13990 3427 13999 3441
rect 13999 3427 14033 3441
rect 14033 3427 14042 3441
rect 14062 3427 14114 3479
rect 13990 3407 13999 3414
rect 13999 3407 14033 3414
rect 14033 3407 14042 3414
rect 13990 3368 14042 3407
rect 13990 3362 13999 3368
rect 13999 3362 14033 3368
rect 14033 3362 14042 3368
rect 14062 3362 14114 3414
rect 13990 3334 13999 3349
rect 13999 3334 14033 3349
rect 14033 3334 14042 3349
rect 13990 3297 14042 3334
rect 14062 3297 14114 3349
rect 13990 3261 13999 3284
rect 13999 3261 14033 3284
rect 14033 3261 14042 3284
rect 13990 3232 14042 3261
rect 14062 3232 14114 3284
rect 13990 3188 13999 3219
rect 13999 3188 14033 3219
rect 14033 3188 14042 3219
rect 13990 3167 14042 3188
rect 14062 3167 14114 3219
rect 13990 3149 14042 3154
rect 13990 3115 13999 3149
rect 13999 3115 14033 3149
rect 14033 3115 14042 3149
rect 13990 3102 14042 3115
rect 14062 3102 14114 3154
rect 13990 3076 14042 3089
rect 13990 3042 13999 3076
rect 13999 3042 14033 3076
rect 14033 3042 14042 3076
rect 13990 3037 14042 3042
rect 14062 3037 14114 3089
rect 13990 3003 14042 3024
rect 13990 2972 13999 3003
rect 13999 2972 14033 3003
rect 14033 2972 14042 3003
rect 14062 2972 14114 3024
rect 14350 2646 14356 2657
rect 14356 2646 14390 2657
rect 14390 2646 14402 2657
rect 14350 2607 14402 2646
rect 14350 2605 14356 2607
rect 14356 2605 14390 2607
rect 14390 2605 14402 2607
rect 14422 2656 14474 2657
rect 14422 2622 14428 2656
rect 14428 2622 14462 2656
rect 14462 2622 14474 2656
rect 14422 2605 14474 2622
rect 14494 2646 14500 2657
rect 14500 2646 14534 2657
rect 14534 2646 14546 2657
rect 14494 2607 14546 2646
rect 14494 2605 14500 2607
rect 14500 2605 14534 2607
rect 14534 2605 14546 2607
rect 14566 2646 14572 2657
rect 14572 2646 14606 2657
rect 14606 2646 14618 2657
rect 14566 2607 14618 2646
rect 14566 2605 14572 2607
rect 14572 2605 14606 2607
rect 14606 2605 14618 2607
rect 14350 2573 14356 2592
rect 14356 2573 14390 2592
rect 14390 2573 14402 2592
rect 14350 2540 14402 2573
rect 14422 2584 14474 2592
rect 14422 2550 14428 2584
rect 14428 2550 14462 2584
rect 14462 2550 14474 2584
rect 14422 2540 14474 2550
rect 14494 2573 14500 2592
rect 14500 2573 14534 2592
rect 14534 2573 14546 2592
rect 14494 2540 14546 2573
rect 14566 2573 14572 2592
rect 14572 2573 14606 2592
rect 14606 2573 14618 2592
rect 14566 2540 14618 2573
rect 14350 2500 14356 2527
rect 14356 2500 14390 2527
rect 14390 2500 14402 2527
rect 14350 2475 14402 2500
rect 14422 2512 14474 2527
rect 14422 2478 14428 2512
rect 14428 2478 14462 2512
rect 14462 2478 14474 2512
rect 14422 2475 14474 2478
rect 14494 2500 14500 2527
rect 14500 2500 14534 2527
rect 14534 2500 14546 2527
rect 14494 2475 14546 2500
rect 14566 2500 14572 2527
rect 14572 2500 14606 2527
rect 14606 2500 14618 2527
rect 14566 2475 14618 2500
rect 14350 2461 14402 2462
rect 14350 2427 14356 2461
rect 14356 2427 14390 2461
rect 14390 2427 14402 2461
rect 14350 2410 14402 2427
rect 14422 2440 14474 2462
rect 14422 2410 14428 2440
rect 14428 2410 14462 2440
rect 14462 2410 14474 2440
rect 14494 2461 14546 2462
rect 14494 2427 14500 2461
rect 14500 2427 14534 2461
rect 14534 2427 14546 2461
rect 14494 2410 14546 2427
rect 14566 2461 14618 2462
rect 14566 2427 14572 2461
rect 14572 2427 14606 2461
rect 14606 2427 14618 2461
rect 14566 2410 14618 2427
rect 14350 2388 14402 2397
rect 14350 2354 14356 2388
rect 14356 2354 14390 2388
rect 14390 2354 14402 2388
rect 14350 2345 14402 2354
rect 14422 2368 14474 2397
rect 14422 2345 14428 2368
rect 14428 2345 14462 2368
rect 14462 2345 14474 2368
rect 14494 2388 14546 2397
rect 14494 2354 14500 2388
rect 14500 2354 14534 2388
rect 14534 2354 14546 2388
rect 14494 2345 14546 2354
rect 14566 2388 14618 2397
rect 14566 2354 14572 2388
rect 14572 2354 14606 2388
rect 14606 2354 14618 2388
rect 14566 2345 14618 2354
rect 14350 2315 14402 2332
rect 14350 2281 14356 2315
rect 14356 2281 14390 2315
rect 14390 2281 14402 2315
rect 14350 2280 14402 2281
rect 14422 2296 14474 2332
rect 14422 2280 14428 2296
rect 14428 2280 14462 2296
rect 14462 2280 14474 2296
rect 14494 2315 14546 2332
rect 14494 2281 14500 2315
rect 14500 2281 14534 2315
rect 14534 2281 14546 2315
rect 14494 2280 14546 2281
rect 14566 2315 14618 2332
rect 14566 2281 14572 2315
rect 14572 2281 14606 2315
rect 14606 2281 14618 2315
rect 14566 2280 14618 2281
rect 14350 2242 14402 2267
rect 14350 2215 14356 2242
rect 14356 2215 14390 2242
rect 14390 2215 14402 2242
rect 14422 2262 14428 2267
rect 14428 2262 14462 2267
rect 14462 2262 14474 2267
rect 14422 2224 14474 2262
rect 14422 2215 14428 2224
rect 14428 2215 14462 2224
rect 14462 2215 14474 2224
rect 14494 2242 14546 2267
rect 14494 2215 14500 2242
rect 14500 2215 14534 2242
rect 14534 2215 14546 2242
rect 14566 2242 14618 2267
rect 14566 2215 14572 2242
rect 14572 2215 14606 2242
rect 14606 2215 14618 2242
rect 14350 2169 14402 2202
rect 14350 2150 14356 2169
rect 14356 2150 14390 2169
rect 14390 2150 14402 2169
rect 14422 2190 14428 2202
rect 14428 2190 14462 2202
rect 14462 2190 14474 2202
rect 14422 2152 14474 2190
rect 14422 2150 14428 2152
rect 14428 2150 14462 2152
rect 14462 2150 14474 2152
rect 14494 2169 14546 2202
rect 14494 2150 14500 2169
rect 14500 2150 14534 2169
rect 14534 2150 14546 2169
rect 14566 2169 14618 2202
rect 14566 2150 14572 2169
rect 14572 2150 14606 2169
rect 14606 2150 14618 2169
rect 14350 2135 14356 2137
rect 14356 2135 14390 2137
rect 14390 2135 14402 2137
rect 14350 2096 14402 2135
rect 14350 2085 14356 2096
rect 14356 2085 14390 2096
rect 14390 2085 14402 2096
rect 14422 2118 14428 2137
rect 14428 2118 14462 2137
rect 14462 2118 14474 2137
rect 14422 2085 14474 2118
rect 14494 2135 14500 2137
rect 14500 2135 14534 2137
rect 14534 2135 14546 2137
rect 14494 2096 14546 2135
rect 14494 2085 14500 2096
rect 14500 2085 14534 2096
rect 14534 2085 14546 2096
rect 14566 2135 14572 2137
rect 14572 2135 14606 2137
rect 14606 2135 14618 2137
rect 14566 2096 14618 2135
rect 14566 2085 14572 2096
rect 14572 2085 14606 2096
rect 14606 2085 14618 2096
rect 14350 2062 14356 2072
rect 14356 2062 14390 2072
rect 14390 2062 14402 2072
rect 14350 2023 14402 2062
rect 14350 2020 14356 2023
rect 14356 2020 14390 2023
rect 14390 2020 14402 2023
rect 14422 2046 14428 2072
rect 14428 2046 14462 2072
rect 14462 2046 14474 2072
rect 14422 2020 14474 2046
rect 14494 2062 14500 2072
rect 14500 2062 14534 2072
rect 14534 2062 14546 2072
rect 14494 2023 14546 2062
rect 14494 2020 14500 2023
rect 14500 2020 14534 2023
rect 14534 2020 14546 2023
rect 14566 2062 14572 2072
rect 14572 2062 14606 2072
rect 14606 2062 14618 2072
rect 14566 2023 14618 2062
rect 14566 2020 14572 2023
rect 14572 2020 14606 2023
rect 14606 2020 14618 2023
rect 14350 1989 14356 2007
rect 14356 1989 14390 2007
rect 14390 1989 14402 2007
rect 14350 1955 14402 1989
rect 14422 1974 14428 2007
rect 14428 1974 14462 2007
rect 14462 1974 14474 2007
rect 14422 1955 14474 1974
rect 14494 1989 14500 2007
rect 14500 1989 14534 2007
rect 14534 1989 14546 2007
rect 14494 1955 14546 1989
rect 14566 1989 14572 2007
rect 14572 1989 14606 2007
rect 14606 1989 14618 2007
rect 14566 1955 14618 1989
rect 14350 1916 14356 1942
rect 14356 1916 14390 1942
rect 14390 1916 14402 1942
rect 14350 1890 14402 1916
rect 14422 1936 14474 1942
rect 14422 1902 14428 1936
rect 14428 1902 14462 1936
rect 14462 1902 14474 1936
rect 14422 1890 14474 1902
rect 14494 1916 14500 1942
rect 14500 1916 14534 1942
rect 14534 1916 14546 1942
rect 14494 1890 14546 1916
rect 14566 1916 14572 1942
rect 14572 1916 14606 1942
rect 14606 1916 14618 1942
rect 14566 1890 14618 1916
rect 14350 1843 14356 1877
rect 14356 1843 14390 1877
rect 14390 1843 14402 1877
rect 14350 1825 14402 1843
rect 14422 1864 14474 1877
rect 14422 1830 14428 1864
rect 14428 1830 14462 1864
rect 14462 1830 14474 1864
rect 14422 1825 14474 1830
rect 14494 1843 14500 1877
rect 14500 1843 14534 1877
rect 14534 1843 14546 1877
rect 14494 1825 14546 1843
rect 14566 1843 14572 1877
rect 14572 1843 14606 1877
rect 14606 1843 14618 1877
rect 14566 1825 14618 1843
rect 14350 1804 14402 1812
rect 14350 1770 14356 1804
rect 14356 1770 14390 1804
rect 14390 1770 14402 1804
rect 14350 1760 14402 1770
rect 14422 1792 14474 1812
rect 14422 1760 14428 1792
rect 14428 1760 14462 1792
rect 14462 1760 14474 1792
rect 14494 1804 14546 1812
rect 14494 1770 14500 1804
rect 14500 1770 14534 1804
rect 14534 1770 14546 1804
rect 14494 1760 14546 1770
rect 14566 1804 14618 1812
rect 14566 1770 14572 1804
rect 14572 1770 14606 1804
rect 14606 1770 14618 1804
rect 14566 1760 14618 1770
rect 14350 1731 14402 1748
rect 14350 1697 14356 1731
rect 14356 1697 14390 1731
rect 14390 1697 14402 1731
rect 14350 1696 14402 1697
rect 14422 1720 14474 1748
rect 14422 1696 14428 1720
rect 14428 1696 14462 1720
rect 14462 1696 14474 1720
rect 14494 1731 14546 1748
rect 14494 1697 14500 1731
rect 14500 1697 14534 1731
rect 14534 1697 14546 1731
rect 14494 1696 14546 1697
rect 14566 1731 14618 1748
rect 14566 1697 14572 1731
rect 14572 1697 14606 1731
rect 14606 1697 14618 1731
rect 14566 1696 14618 1697
rect 14350 1657 14402 1684
rect 14350 1632 14356 1657
rect 14356 1632 14390 1657
rect 14390 1632 14402 1657
rect 14422 1648 14474 1684
rect 14422 1632 14428 1648
rect 14428 1632 14462 1648
rect 14462 1632 14474 1648
rect 14494 1658 14546 1684
rect 14494 1632 14500 1658
rect 14500 1632 14534 1658
rect 14534 1632 14546 1658
rect 14566 1658 14618 1684
rect 14566 1632 14572 1658
rect 14572 1632 14606 1658
rect 14606 1632 14618 1658
rect 14350 1583 14402 1620
rect 14350 1568 14356 1583
rect 14356 1568 14390 1583
rect 14390 1568 14402 1583
rect 14422 1614 14428 1620
rect 14428 1614 14462 1620
rect 14462 1614 14474 1620
rect 14422 1576 14474 1614
rect 14422 1568 14428 1576
rect 14428 1568 14462 1576
rect 14462 1568 14474 1576
rect 14494 1585 14546 1620
rect 14494 1568 14500 1585
rect 14500 1568 14534 1585
rect 14534 1568 14546 1585
rect 14566 1585 14618 1620
rect 14566 1568 14572 1585
rect 14572 1568 14606 1585
rect 14606 1568 14618 1585
<< metal2 >>
rect 1061 4119 14114 4125
rect 1061 4067 1066 4119
rect 1118 4067 1130 4119
rect 1182 4067 1194 4119
rect 1246 4067 2058 4119
rect 2110 4067 2122 4119
rect 2174 4067 2186 4119
rect 2238 4067 3050 4119
rect 3102 4067 3114 4119
rect 3166 4067 3178 4119
rect 3230 4067 4042 4119
rect 4094 4067 4106 4119
rect 4158 4067 4170 4119
rect 4222 4067 5034 4119
rect 5086 4067 5098 4119
rect 5150 4067 5162 4119
rect 5214 4067 6026 4119
rect 6078 4067 6090 4119
rect 6142 4067 6154 4119
rect 6206 4067 7018 4119
rect 7070 4067 7082 4119
rect 7134 4067 7146 4119
rect 7198 4067 8010 4119
rect 8062 4067 8074 4119
rect 8126 4067 8138 4119
rect 8190 4067 9002 4119
rect 9054 4067 9066 4119
rect 9118 4067 9130 4119
rect 9182 4067 9994 4119
rect 10046 4067 10058 4119
rect 10110 4067 10122 4119
rect 10174 4067 10986 4119
rect 11038 4067 11050 4119
rect 11102 4067 11114 4119
rect 11166 4067 11978 4119
rect 12030 4067 12042 4119
rect 12094 4067 12106 4119
rect 12158 4067 12970 4119
rect 13022 4067 13034 4119
rect 13086 4067 13098 4119
rect 13150 4067 13990 4119
rect 14042 4067 14062 4119
rect 1061 4055 14114 4067
rect 1061 4054 13990 4055
rect 1061 4002 1066 4054
rect 1118 4002 1130 4054
rect 1182 4002 1194 4054
rect 1246 4002 2058 4054
rect 2110 4002 2122 4054
rect 2174 4002 2186 4054
rect 2238 4002 3050 4054
rect 3102 4002 3114 4054
rect 3166 4002 3178 4054
rect 3230 4002 4042 4054
rect 4094 4002 4106 4054
rect 4158 4002 4170 4054
rect 4222 4002 5034 4054
rect 5086 4002 5098 4054
rect 5150 4002 5162 4054
rect 5214 4002 6026 4054
rect 6078 4002 6090 4054
rect 6142 4002 6154 4054
rect 6206 4002 7018 4054
rect 7070 4002 7082 4054
rect 7134 4002 7146 4054
rect 7198 4002 8010 4054
rect 8062 4002 8074 4054
rect 8126 4002 8138 4054
rect 8190 4002 9002 4054
rect 9054 4002 9066 4054
rect 9118 4002 9130 4054
rect 9182 4002 9994 4054
rect 10046 4002 10058 4054
rect 10110 4002 10122 4054
rect 10174 4002 10986 4054
rect 11038 4002 11050 4054
rect 11102 4002 11114 4054
rect 11166 4002 11978 4054
rect 12030 4002 12042 4054
rect 12094 4002 12106 4054
rect 12158 4002 12970 4054
rect 13022 4002 13034 4054
rect 13086 4002 13098 4054
rect 13150 4003 13990 4054
rect 14042 4003 14062 4055
rect 13150 4002 14114 4003
rect 1061 3991 14114 4002
rect 1061 3989 13990 3991
rect 1061 3937 1066 3989
rect 1118 3937 1130 3989
rect 1182 3937 1194 3989
rect 1246 3937 2058 3989
rect 2110 3937 2122 3989
rect 2174 3937 2186 3989
rect 2238 3937 3050 3989
rect 3102 3937 3114 3989
rect 3166 3937 3178 3989
rect 3230 3937 4042 3989
rect 4094 3937 4106 3989
rect 4158 3937 4170 3989
rect 4222 3937 5034 3989
rect 5086 3937 5098 3989
rect 5150 3937 5162 3989
rect 5214 3937 6026 3989
rect 6078 3937 6090 3989
rect 6142 3937 6154 3989
rect 6206 3937 7018 3989
rect 7070 3937 7082 3989
rect 7134 3937 7146 3989
rect 7198 3937 8010 3989
rect 8062 3937 8074 3989
rect 8126 3937 8138 3989
rect 8190 3937 9002 3989
rect 9054 3937 9066 3989
rect 9118 3937 9130 3989
rect 9182 3937 9994 3989
rect 10046 3937 10058 3989
rect 10110 3937 10122 3989
rect 10174 3937 10986 3989
rect 11038 3937 11050 3989
rect 11102 3937 11114 3989
rect 11166 3937 11978 3989
rect 12030 3937 12042 3989
rect 12094 3937 12106 3989
rect 12158 3937 12970 3989
rect 13022 3937 13034 3989
rect 13086 3937 13098 3989
rect 13150 3939 13990 3989
rect 14042 3939 14062 3991
rect 13150 3937 14114 3939
rect 1061 3927 14114 3937
rect 1061 3924 13990 3927
rect 1061 3872 1066 3924
rect 1118 3872 1130 3924
rect 1182 3872 1194 3924
rect 1246 3872 2058 3924
rect 2110 3872 2122 3924
rect 2174 3872 2186 3924
rect 2238 3872 3050 3924
rect 3102 3872 3114 3924
rect 3166 3872 3178 3924
rect 3230 3872 4042 3924
rect 4094 3872 4106 3924
rect 4158 3872 4170 3924
rect 4222 3872 5034 3924
rect 5086 3872 5098 3924
rect 5150 3872 5162 3924
rect 5214 3872 6026 3924
rect 6078 3872 6090 3924
rect 6142 3872 6154 3924
rect 6206 3872 7018 3924
rect 7070 3872 7082 3924
rect 7134 3872 7146 3924
rect 7198 3872 8010 3924
rect 8062 3872 8074 3924
rect 8126 3872 8138 3924
rect 8190 3872 9002 3924
rect 9054 3872 9066 3924
rect 9118 3872 9130 3924
rect 9182 3872 9994 3924
rect 10046 3872 10058 3924
rect 10110 3872 10122 3924
rect 10174 3872 10986 3924
rect 11038 3872 11050 3924
rect 11102 3872 11114 3924
rect 11166 3872 11978 3924
rect 12030 3872 12042 3924
rect 12094 3872 12106 3924
rect 12158 3872 12970 3924
rect 13022 3872 13034 3924
rect 13086 3872 13098 3924
rect 13150 3875 13990 3924
rect 14042 3875 14062 3927
rect 13150 3872 14114 3875
rect 1061 3863 14114 3872
rect 1061 3859 13990 3863
rect 1061 3807 1066 3859
rect 1118 3807 1130 3859
rect 1182 3807 1194 3859
rect 1246 3807 2058 3859
rect 2110 3807 2122 3859
rect 2174 3807 2186 3859
rect 2238 3807 3050 3859
rect 3102 3807 3114 3859
rect 3166 3807 3178 3859
rect 3230 3807 4042 3859
rect 4094 3807 4106 3859
rect 4158 3807 4170 3859
rect 4222 3807 5034 3859
rect 5086 3807 5098 3859
rect 5150 3807 5162 3859
rect 5214 3807 6026 3859
rect 6078 3807 6090 3859
rect 6142 3807 6154 3859
rect 6206 3807 7018 3859
rect 7070 3807 7082 3859
rect 7134 3807 7146 3859
rect 7198 3807 8010 3859
rect 8062 3807 8074 3859
rect 8126 3807 8138 3859
rect 8190 3807 9002 3859
rect 9054 3807 9066 3859
rect 9118 3807 9130 3859
rect 9182 3807 9994 3859
rect 10046 3807 10058 3859
rect 10110 3807 10122 3859
rect 10174 3807 10986 3859
rect 11038 3807 11050 3859
rect 11102 3807 11114 3859
rect 11166 3807 11978 3859
rect 12030 3807 12042 3859
rect 12094 3807 12106 3859
rect 12158 3807 12970 3859
rect 13022 3807 13034 3859
rect 13086 3807 13098 3859
rect 13150 3811 13990 3859
rect 14042 3811 14062 3863
rect 13150 3807 14114 3811
rect 1061 3799 14114 3807
rect 1061 3794 13990 3799
rect 1061 3742 1066 3794
rect 1118 3742 1130 3794
rect 1182 3742 1194 3794
rect 1246 3742 2058 3794
rect 2110 3742 2122 3794
rect 2174 3742 2186 3794
rect 2238 3742 3050 3794
rect 3102 3742 3114 3794
rect 3166 3742 3178 3794
rect 3230 3742 4042 3794
rect 4094 3742 4106 3794
rect 4158 3742 4170 3794
rect 4222 3742 5034 3794
rect 5086 3742 5098 3794
rect 5150 3742 5162 3794
rect 5214 3742 6026 3794
rect 6078 3742 6090 3794
rect 6142 3742 6154 3794
rect 6206 3742 7018 3794
rect 7070 3742 7082 3794
rect 7134 3742 7146 3794
rect 7198 3742 8010 3794
rect 8062 3742 8074 3794
rect 8126 3742 8138 3794
rect 8190 3742 9002 3794
rect 9054 3742 9066 3794
rect 9118 3742 9130 3794
rect 9182 3742 9994 3794
rect 10046 3742 10058 3794
rect 10110 3742 10122 3794
rect 10174 3742 10986 3794
rect 11038 3742 11050 3794
rect 11102 3742 11114 3794
rect 11166 3742 11978 3794
rect 12030 3742 12042 3794
rect 12094 3742 12106 3794
rect 12158 3742 12970 3794
rect 13022 3742 13034 3794
rect 13086 3742 13098 3794
rect 13150 3747 13990 3794
rect 14042 3747 14062 3799
rect 13150 3742 14114 3747
rect 1061 3735 14114 3742
rect 1061 3729 13990 3735
rect 1061 3677 1066 3729
rect 1118 3677 1130 3729
rect 1182 3677 1194 3729
rect 1246 3677 2058 3729
rect 2110 3677 2122 3729
rect 2174 3677 2186 3729
rect 2238 3677 3050 3729
rect 3102 3677 3114 3729
rect 3166 3677 3178 3729
rect 3230 3677 4042 3729
rect 4094 3677 4106 3729
rect 4158 3677 4170 3729
rect 4222 3677 5034 3729
rect 5086 3677 5098 3729
rect 5150 3677 5162 3729
rect 5214 3677 6026 3729
rect 6078 3677 6090 3729
rect 6142 3677 6154 3729
rect 6206 3677 7018 3729
rect 7070 3677 7082 3729
rect 7134 3677 7146 3729
rect 7198 3677 8010 3729
rect 8062 3677 8074 3729
rect 8126 3677 8138 3729
rect 8190 3677 9002 3729
rect 9054 3677 9066 3729
rect 9118 3677 9130 3729
rect 9182 3677 9994 3729
rect 10046 3677 10058 3729
rect 10110 3677 10122 3729
rect 10174 3677 10986 3729
rect 11038 3677 11050 3729
rect 11102 3677 11114 3729
rect 11166 3677 11978 3729
rect 12030 3677 12042 3729
rect 12094 3677 12106 3729
rect 12158 3677 12970 3729
rect 13022 3677 13034 3729
rect 13086 3677 13098 3729
rect 13150 3683 13990 3729
rect 14042 3683 14062 3735
rect 13150 3677 14114 3683
rect 1061 3671 14114 3677
rect 1061 3664 13990 3671
rect 1061 2972 1066 3664
rect 1246 2972 2058 3664
rect 2238 2972 3050 3664
rect 3230 2972 4042 3664
rect 4222 2972 5034 3664
rect 5214 2972 6026 3664
rect 6206 2972 7018 3664
rect 7198 2972 8010 3664
rect 8190 2972 9002 3664
rect 9182 2972 9994 3664
rect 10174 2972 10986 3664
rect 11166 2972 11978 3664
rect 12158 2972 12970 3664
rect 13150 3619 13990 3664
rect 14042 3619 14062 3671
rect 13150 3607 14114 3619
rect 13150 3555 13990 3607
rect 14042 3555 14062 3607
rect 13150 3543 14114 3555
rect 13150 3491 13990 3543
rect 14042 3491 14062 3543
rect 13150 3479 14114 3491
rect 13150 3427 13990 3479
rect 14042 3427 14062 3479
rect 13150 3414 14114 3427
rect 13150 3362 13990 3414
rect 14042 3362 14062 3414
rect 13150 3349 14114 3362
rect 13150 3297 13990 3349
rect 14042 3297 14062 3349
rect 13150 3284 14114 3297
rect 13150 3232 13990 3284
rect 14042 3232 14062 3284
rect 13150 3219 14114 3232
rect 13150 3167 13990 3219
rect 14042 3167 14062 3219
rect 13150 3154 14114 3167
rect 13150 3102 13990 3154
rect 14042 3102 14062 3154
rect 13150 3089 14114 3102
rect 13150 3037 13990 3089
rect 14042 3037 14062 3089
rect 13150 3024 14114 3037
rect 13150 2972 13990 3024
rect 14042 2972 14062 3024
rect 1061 2966 14114 2972
rect 558 2657 14618 2663
rect 610 2605 646 2657
rect 698 2605 734 2657
rect 786 2605 1562 2657
rect 1614 2605 1626 2657
rect 1678 2605 1690 2657
rect 1742 2605 2554 2657
rect 2606 2605 2618 2657
rect 2670 2605 2682 2657
rect 2734 2605 3546 2657
rect 3598 2605 3610 2657
rect 3662 2605 3674 2657
rect 3726 2605 4538 2657
rect 4590 2605 4602 2657
rect 4654 2605 4666 2657
rect 4718 2605 5530 2657
rect 5582 2605 5594 2657
rect 5646 2605 5658 2657
rect 5710 2605 6522 2657
rect 6574 2605 6586 2657
rect 6638 2605 6650 2657
rect 6702 2605 7514 2657
rect 7566 2605 7578 2657
rect 7630 2605 7642 2657
rect 7694 2605 8506 2657
rect 8558 2605 8570 2657
rect 8622 2605 8634 2657
rect 8686 2605 9498 2657
rect 9550 2605 9562 2657
rect 9614 2605 9626 2657
rect 9678 2605 10490 2657
rect 10542 2605 10554 2657
rect 10606 2605 10618 2657
rect 10670 2605 11482 2657
rect 11534 2605 11546 2657
rect 11598 2605 11610 2657
rect 11662 2605 12474 2657
rect 12526 2605 12538 2657
rect 12590 2605 12602 2657
rect 12654 2605 13466 2657
rect 13518 2605 13530 2657
rect 13582 2605 13594 2657
rect 13646 2605 14350 2657
rect 14402 2605 14422 2657
rect 14474 2605 14494 2657
rect 14546 2605 14566 2657
rect 558 2592 14618 2605
rect 610 2540 646 2592
rect 698 2540 734 2592
rect 786 2540 1562 2592
rect 1614 2540 1626 2592
rect 1678 2540 1690 2592
rect 1742 2540 2554 2592
rect 2606 2540 2618 2592
rect 2670 2540 2682 2592
rect 2734 2540 3546 2592
rect 3598 2540 3610 2592
rect 3662 2540 3674 2592
rect 3726 2540 4538 2592
rect 4590 2540 4602 2592
rect 4654 2540 4666 2592
rect 4718 2540 5530 2592
rect 5582 2540 5594 2592
rect 5646 2540 5658 2592
rect 5710 2540 6522 2592
rect 6574 2540 6586 2592
rect 6638 2540 6650 2592
rect 6702 2540 7514 2592
rect 7566 2540 7578 2592
rect 7630 2540 7642 2592
rect 7694 2540 8506 2592
rect 8558 2540 8570 2592
rect 8622 2540 8634 2592
rect 8686 2540 9498 2592
rect 9550 2540 9562 2592
rect 9614 2540 9626 2592
rect 9678 2540 10490 2592
rect 10542 2540 10554 2592
rect 10606 2540 10618 2592
rect 10670 2540 11482 2592
rect 11534 2540 11546 2592
rect 11598 2540 11610 2592
rect 11662 2540 12474 2592
rect 12526 2540 12538 2592
rect 12590 2540 12602 2592
rect 12654 2540 13466 2592
rect 13518 2540 13530 2592
rect 13582 2540 13594 2592
rect 13646 2540 14350 2592
rect 14402 2540 14422 2592
rect 14474 2540 14494 2592
rect 14546 2540 14566 2592
rect 558 2527 14618 2540
rect 610 2475 646 2527
rect 698 2475 734 2527
rect 786 2475 1562 2527
rect 1614 2475 1626 2527
rect 1678 2475 1690 2527
rect 1742 2475 2554 2527
rect 2606 2475 2618 2527
rect 2670 2475 2682 2527
rect 2734 2475 3546 2527
rect 3598 2475 3610 2527
rect 3662 2475 3674 2527
rect 3726 2475 4538 2527
rect 4590 2475 4602 2527
rect 4654 2475 4666 2527
rect 4718 2475 5530 2527
rect 5582 2475 5594 2527
rect 5646 2475 5658 2527
rect 5710 2475 6522 2527
rect 6574 2475 6586 2527
rect 6638 2475 6650 2527
rect 6702 2475 7514 2527
rect 7566 2475 7578 2527
rect 7630 2475 7642 2527
rect 7694 2475 8506 2527
rect 8558 2475 8570 2527
rect 8622 2475 8634 2527
rect 8686 2475 9498 2527
rect 9550 2475 9562 2527
rect 9614 2475 9626 2527
rect 9678 2475 10490 2527
rect 10542 2475 10554 2527
rect 10606 2475 10618 2527
rect 10670 2475 11482 2527
rect 11534 2475 11546 2527
rect 11598 2475 11610 2527
rect 11662 2475 12474 2527
rect 12526 2475 12538 2527
rect 12590 2475 12602 2527
rect 12654 2475 13466 2527
rect 13518 2475 13530 2527
rect 13582 2475 13594 2527
rect 13646 2475 14350 2527
rect 14402 2475 14422 2527
rect 14474 2475 14494 2527
rect 14546 2475 14566 2527
rect 558 2462 14618 2475
rect 610 2410 646 2462
rect 698 2410 734 2462
rect 786 2410 1562 2462
rect 1614 2410 1626 2462
rect 1678 2410 1690 2462
rect 1742 2410 2554 2462
rect 2606 2410 2618 2462
rect 2670 2410 2682 2462
rect 2734 2410 3546 2462
rect 3598 2410 3610 2462
rect 3662 2410 3674 2462
rect 3726 2410 4538 2462
rect 4590 2410 4602 2462
rect 4654 2410 4666 2462
rect 4718 2410 5530 2462
rect 5582 2410 5594 2462
rect 5646 2410 5658 2462
rect 5710 2410 6522 2462
rect 6574 2410 6586 2462
rect 6638 2410 6650 2462
rect 6702 2410 7514 2462
rect 7566 2410 7578 2462
rect 7630 2410 7642 2462
rect 7694 2410 8506 2462
rect 8558 2410 8570 2462
rect 8622 2410 8634 2462
rect 8686 2410 9498 2462
rect 9550 2410 9562 2462
rect 9614 2410 9626 2462
rect 9678 2410 10490 2462
rect 10542 2410 10554 2462
rect 10606 2410 10618 2462
rect 10670 2410 11482 2462
rect 11534 2410 11546 2462
rect 11598 2410 11610 2462
rect 11662 2410 12474 2462
rect 12526 2410 12538 2462
rect 12590 2410 12602 2462
rect 12654 2410 13466 2462
rect 13518 2410 13530 2462
rect 13582 2410 13594 2462
rect 13646 2410 14350 2462
rect 14402 2410 14422 2462
rect 14474 2410 14494 2462
rect 14546 2410 14566 2462
rect 558 2397 14618 2410
rect 610 2345 646 2397
rect 698 2345 734 2397
rect 786 2345 1562 2397
rect 1614 2345 1626 2397
rect 1678 2345 1690 2397
rect 1742 2345 2554 2397
rect 2606 2345 2618 2397
rect 2670 2345 2682 2397
rect 2734 2345 3546 2397
rect 3598 2345 3610 2397
rect 3662 2345 3674 2397
rect 3726 2345 4538 2397
rect 4590 2345 4602 2397
rect 4654 2345 4666 2397
rect 4718 2345 5530 2397
rect 5582 2345 5594 2397
rect 5646 2345 5658 2397
rect 5710 2345 6522 2397
rect 6574 2345 6586 2397
rect 6638 2345 6650 2397
rect 6702 2345 7514 2397
rect 7566 2345 7578 2397
rect 7630 2345 7642 2397
rect 7694 2345 8506 2397
rect 8558 2345 8570 2397
rect 8622 2345 8634 2397
rect 8686 2345 9498 2397
rect 9550 2345 9562 2397
rect 9614 2345 9626 2397
rect 9678 2345 10490 2397
rect 10542 2345 10554 2397
rect 10606 2345 10618 2397
rect 10670 2345 11482 2397
rect 11534 2345 11546 2397
rect 11598 2345 11610 2397
rect 11662 2345 12474 2397
rect 12526 2345 12538 2397
rect 12590 2345 12602 2397
rect 12654 2345 13466 2397
rect 13518 2345 13530 2397
rect 13582 2345 13594 2397
rect 13646 2345 14350 2397
rect 14402 2345 14422 2397
rect 14474 2345 14494 2397
rect 14546 2345 14566 2397
rect 558 2332 14618 2345
rect 610 2280 646 2332
rect 698 2280 734 2332
rect 786 2280 1562 2332
rect 1614 2280 1626 2332
rect 1678 2280 1690 2332
rect 1742 2280 2554 2332
rect 2606 2280 2618 2332
rect 2670 2280 2682 2332
rect 2734 2280 3546 2332
rect 3598 2280 3610 2332
rect 3662 2280 3674 2332
rect 3726 2280 4538 2332
rect 4590 2280 4602 2332
rect 4654 2280 4666 2332
rect 4718 2280 5530 2332
rect 5582 2280 5594 2332
rect 5646 2280 5658 2332
rect 5710 2280 6522 2332
rect 6574 2280 6586 2332
rect 6638 2280 6650 2332
rect 6702 2280 7514 2332
rect 7566 2280 7578 2332
rect 7630 2280 7642 2332
rect 7694 2280 8506 2332
rect 8558 2280 8570 2332
rect 8622 2280 8634 2332
rect 8686 2280 9498 2332
rect 9550 2280 9562 2332
rect 9614 2280 9626 2332
rect 9678 2280 10490 2332
rect 10542 2280 10554 2332
rect 10606 2280 10618 2332
rect 10670 2280 11482 2332
rect 11534 2280 11546 2332
rect 11598 2280 11610 2332
rect 11662 2280 12474 2332
rect 12526 2280 12538 2332
rect 12590 2280 12602 2332
rect 12654 2280 13466 2332
rect 13518 2280 13530 2332
rect 13582 2280 13594 2332
rect 13646 2280 14350 2332
rect 14402 2280 14422 2332
rect 14474 2280 14494 2332
rect 14546 2280 14566 2332
rect 558 2267 14618 2280
rect 610 2215 646 2267
rect 698 2215 734 2267
rect 786 2215 1562 2267
rect 1614 2215 1626 2267
rect 1678 2215 1690 2267
rect 1742 2215 2554 2267
rect 2606 2215 2618 2267
rect 2670 2215 2682 2267
rect 2734 2215 3546 2267
rect 3598 2215 3610 2267
rect 3662 2215 3674 2267
rect 3726 2215 4538 2267
rect 4590 2215 4602 2267
rect 4654 2215 4666 2267
rect 4718 2215 5530 2267
rect 5582 2215 5594 2267
rect 5646 2215 5658 2267
rect 5710 2215 6522 2267
rect 6574 2215 6586 2267
rect 6638 2215 6650 2267
rect 6702 2215 7514 2267
rect 7566 2215 7578 2267
rect 7630 2215 7642 2267
rect 7694 2215 8506 2267
rect 8558 2215 8570 2267
rect 8622 2215 8634 2267
rect 8686 2215 9498 2267
rect 9550 2215 9562 2267
rect 9614 2215 9626 2267
rect 9678 2215 10490 2267
rect 10542 2215 10554 2267
rect 10606 2215 10618 2267
rect 10670 2215 11482 2267
rect 11534 2215 11546 2267
rect 11598 2215 11610 2267
rect 11662 2215 12474 2267
rect 12526 2215 12538 2267
rect 12590 2215 12602 2267
rect 12654 2215 13466 2267
rect 13518 2215 13530 2267
rect 13582 2215 13594 2267
rect 13646 2215 14350 2267
rect 14402 2215 14422 2267
rect 14474 2215 14494 2267
rect 14546 2215 14566 2267
rect 558 2202 14618 2215
rect 610 2150 646 2202
rect 698 2150 734 2202
rect 786 2150 1562 2202
rect 1614 2150 1626 2202
rect 1678 2150 1690 2202
rect 1742 2150 2554 2202
rect 2606 2150 2618 2202
rect 2670 2150 2682 2202
rect 2734 2150 3546 2202
rect 3598 2150 3610 2202
rect 3662 2150 3674 2202
rect 3726 2150 4538 2202
rect 4590 2150 4602 2202
rect 4654 2150 4666 2202
rect 4718 2150 5530 2202
rect 5582 2150 5594 2202
rect 5646 2150 5658 2202
rect 5710 2150 6522 2202
rect 6574 2150 6586 2202
rect 6638 2150 6650 2202
rect 6702 2150 7514 2202
rect 7566 2150 7578 2202
rect 7630 2150 7642 2202
rect 7694 2150 8506 2202
rect 8558 2150 8570 2202
rect 8622 2150 8634 2202
rect 8686 2150 9498 2202
rect 9550 2150 9562 2202
rect 9614 2150 9626 2202
rect 9678 2150 10490 2202
rect 10542 2150 10554 2202
rect 10606 2150 10618 2202
rect 10670 2150 11482 2202
rect 11534 2150 11546 2202
rect 11598 2150 11610 2202
rect 11662 2150 12474 2202
rect 12526 2150 12538 2202
rect 12590 2150 12602 2202
rect 12654 2150 13466 2202
rect 13518 2150 13530 2202
rect 13582 2150 13594 2202
rect 13646 2150 14350 2202
rect 14402 2150 14422 2202
rect 14474 2150 14494 2202
rect 14546 2150 14566 2202
rect 558 2137 14618 2150
rect 610 2085 646 2137
rect 698 2085 734 2137
rect 786 2085 1562 2137
rect 1614 2085 1626 2137
rect 1678 2085 1690 2137
rect 1742 2085 2554 2137
rect 2606 2085 2618 2137
rect 2670 2085 2682 2137
rect 2734 2085 3546 2137
rect 3598 2085 3610 2137
rect 3662 2085 3674 2137
rect 3726 2085 4538 2137
rect 4590 2085 4602 2137
rect 4654 2085 4666 2137
rect 4718 2085 5530 2137
rect 5582 2085 5594 2137
rect 5646 2085 5658 2137
rect 5710 2085 6522 2137
rect 6574 2085 6586 2137
rect 6638 2085 6650 2137
rect 6702 2085 7514 2137
rect 7566 2085 7578 2137
rect 7630 2085 7642 2137
rect 7694 2085 8506 2137
rect 8558 2085 8570 2137
rect 8622 2085 8634 2137
rect 8686 2085 9498 2137
rect 9550 2085 9562 2137
rect 9614 2085 9626 2137
rect 9678 2085 10490 2137
rect 10542 2085 10554 2137
rect 10606 2085 10618 2137
rect 10670 2085 11482 2137
rect 11534 2085 11546 2137
rect 11598 2085 11610 2137
rect 11662 2085 12474 2137
rect 12526 2085 12538 2137
rect 12590 2085 12602 2137
rect 12654 2085 13466 2137
rect 13518 2085 13530 2137
rect 13582 2085 13594 2137
rect 13646 2085 14350 2137
rect 14402 2085 14422 2137
rect 14474 2085 14494 2137
rect 14546 2085 14566 2137
rect 558 2072 14618 2085
rect 610 2020 646 2072
rect 698 2020 734 2072
rect 786 2020 1562 2072
rect 1614 2020 1626 2072
rect 1678 2020 1690 2072
rect 1742 2020 2554 2072
rect 2606 2020 2618 2072
rect 2670 2020 2682 2072
rect 2734 2020 3546 2072
rect 3598 2020 3610 2072
rect 3662 2020 3674 2072
rect 3726 2020 4538 2072
rect 4590 2020 4602 2072
rect 4654 2020 4666 2072
rect 4718 2020 5530 2072
rect 5582 2020 5594 2072
rect 5646 2020 5658 2072
rect 5710 2020 6522 2072
rect 6574 2020 6586 2072
rect 6638 2020 6650 2072
rect 6702 2020 7514 2072
rect 7566 2020 7578 2072
rect 7630 2020 7642 2072
rect 7694 2020 8506 2072
rect 8558 2020 8570 2072
rect 8622 2020 8634 2072
rect 8686 2020 9498 2072
rect 9550 2020 9562 2072
rect 9614 2020 9626 2072
rect 9678 2020 10490 2072
rect 10542 2020 10554 2072
rect 10606 2020 10618 2072
rect 10670 2020 11482 2072
rect 11534 2020 11546 2072
rect 11598 2020 11610 2072
rect 11662 2020 12474 2072
rect 12526 2020 12538 2072
rect 12590 2020 12602 2072
rect 12654 2020 13466 2072
rect 13518 2020 13530 2072
rect 13582 2020 13594 2072
rect 13646 2020 14350 2072
rect 14402 2020 14422 2072
rect 14474 2020 14494 2072
rect 14546 2020 14566 2072
rect 558 2007 14618 2020
rect 610 1955 646 2007
rect 698 1955 734 2007
rect 786 1955 1562 2007
rect 1614 1955 1626 2007
rect 1678 1955 1690 2007
rect 1742 1955 2554 2007
rect 2606 1955 2618 2007
rect 2670 1955 2682 2007
rect 2734 1955 3546 2007
rect 3598 1955 3610 2007
rect 3662 1955 3674 2007
rect 3726 1955 4538 2007
rect 4590 1955 4602 2007
rect 4654 1955 4666 2007
rect 4718 1955 5530 2007
rect 5582 1955 5594 2007
rect 5646 1955 5658 2007
rect 5710 1955 6522 2007
rect 6574 1955 6586 2007
rect 6638 1955 6650 2007
rect 6702 1955 7514 2007
rect 7566 1955 7578 2007
rect 7630 1955 7642 2007
rect 7694 1955 8506 2007
rect 8558 1955 8570 2007
rect 8622 1955 8634 2007
rect 8686 1955 9498 2007
rect 9550 1955 9562 2007
rect 9614 1955 9626 2007
rect 9678 1955 10490 2007
rect 10542 1955 10554 2007
rect 10606 1955 10618 2007
rect 10670 1955 11482 2007
rect 11534 1955 11546 2007
rect 11598 1955 11610 2007
rect 11662 1955 12474 2007
rect 12526 1955 12538 2007
rect 12590 1955 12602 2007
rect 12654 1955 13466 2007
rect 13518 1955 13530 2007
rect 13582 1955 13594 2007
rect 13646 1955 14350 2007
rect 14402 1955 14422 2007
rect 14474 1955 14494 2007
rect 14546 1955 14566 2007
rect 558 1942 14618 1955
rect 610 1890 646 1942
rect 698 1890 734 1942
rect 786 1890 1562 1942
rect 1614 1890 1626 1942
rect 1678 1890 1690 1942
rect 1742 1890 2554 1942
rect 2606 1890 2618 1942
rect 2670 1890 2682 1942
rect 2734 1890 3546 1942
rect 3598 1890 3610 1942
rect 3662 1890 3674 1942
rect 3726 1890 4538 1942
rect 4590 1890 4602 1942
rect 4654 1890 4666 1942
rect 4718 1890 5530 1942
rect 5582 1890 5594 1942
rect 5646 1890 5658 1942
rect 5710 1890 6522 1942
rect 6574 1890 6586 1942
rect 6638 1890 6650 1942
rect 6702 1890 7514 1942
rect 7566 1890 7578 1942
rect 7630 1890 7642 1942
rect 7694 1890 8506 1942
rect 8558 1890 8570 1942
rect 8622 1890 8634 1942
rect 8686 1890 9498 1942
rect 9550 1890 9562 1942
rect 9614 1890 9626 1942
rect 9678 1890 10490 1942
rect 10542 1890 10554 1942
rect 10606 1890 10618 1942
rect 10670 1890 11482 1942
rect 11534 1890 11546 1942
rect 11598 1890 11610 1942
rect 11662 1890 12474 1942
rect 12526 1890 12538 1942
rect 12590 1890 12602 1942
rect 12654 1890 13466 1942
rect 13518 1890 13530 1942
rect 13582 1890 13594 1942
rect 13646 1890 14350 1942
rect 14402 1890 14422 1942
rect 14474 1890 14494 1942
rect 14546 1890 14566 1942
rect 558 1877 14618 1890
rect 610 1825 646 1877
rect 698 1825 734 1877
rect 786 1825 1562 1877
rect 1614 1825 1626 1877
rect 1678 1825 1690 1877
rect 1742 1825 2554 1877
rect 2606 1825 2618 1877
rect 2670 1825 2682 1877
rect 2734 1825 3546 1877
rect 3598 1825 3610 1877
rect 3662 1825 3674 1877
rect 3726 1825 4538 1877
rect 4590 1825 4602 1877
rect 4654 1825 4666 1877
rect 4718 1825 5530 1877
rect 5582 1825 5594 1877
rect 5646 1825 5658 1877
rect 5710 1825 6522 1877
rect 6574 1825 6586 1877
rect 6638 1825 6650 1877
rect 6702 1825 7514 1877
rect 7566 1825 7578 1877
rect 7630 1825 7642 1877
rect 7694 1825 8506 1877
rect 8558 1825 8570 1877
rect 8622 1825 8634 1877
rect 8686 1825 9498 1877
rect 9550 1825 9562 1877
rect 9614 1825 9626 1877
rect 9678 1825 10490 1877
rect 10542 1825 10554 1877
rect 10606 1825 10618 1877
rect 10670 1825 11482 1877
rect 11534 1825 11546 1877
rect 11598 1825 11610 1877
rect 11662 1825 12474 1877
rect 12526 1825 12538 1877
rect 12590 1825 12602 1877
rect 12654 1825 13466 1877
rect 13518 1825 13530 1877
rect 13582 1825 13594 1877
rect 13646 1825 14350 1877
rect 14402 1825 14422 1877
rect 14474 1825 14494 1877
rect 14546 1825 14566 1877
rect 558 1812 14618 1825
rect 610 1760 646 1812
rect 698 1760 734 1812
rect 786 1760 1562 1812
rect 558 1748 1562 1760
rect 610 1696 646 1748
rect 698 1696 734 1748
rect 786 1696 1562 1748
rect 558 1684 1562 1696
rect 610 1632 646 1684
rect 698 1632 734 1684
rect 786 1632 1562 1684
rect 558 1620 1562 1632
rect 610 1568 646 1620
rect 698 1568 734 1620
rect 786 1568 1562 1620
rect 1742 1568 2554 1812
rect 2734 1568 3546 1812
rect 3726 1568 4538 1812
rect 4718 1568 5530 1812
rect 5710 1568 6522 1812
rect 6702 1568 7514 1812
rect 7694 1568 8506 1812
rect 8686 1568 9498 1812
rect 9678 1568 10490 1812
rect 10670 1568 11482 1812
rect 11662 1568 12474 1812
rect 12654 1568 13466 1812
rect 13646 1760 14350 1812
rect 14402 1760 14422 1812
rect 14474 1760 14494 1812
rect 14546 1760 14566 1812
rect 13646 1748 14618 1760
rect 13646 1696 14350 1748
rect 14402 1696 14422 1748
rect 14474 1696 14494 1748
rect 14546 1696 14566 1748
rect 13646 1684 14618 1696
rect 13646 1632 14350 1684
rect 14402 1632 14422 1684
rect 14474 1632 14494 1684
rect 14546 1632 14566 1684
rect 13646 1620 14618 1632
rect 13646 1568 14350 1620
rect 14402 1568 14422 1620
rect 14474 1568 14494 1620
rect 14546 1568 14566 1620
rect 558 1562 14618 1568
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_0
timestamp 1681267127
transform -1 0 8164 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_1
timestamp 1681267127
transform 1 0 8036 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_2
timestamp 1681267127
transform -1 0 7172 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_3
timestamp 1681267127
transform -1 0 6180 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_4
timestamp 1681267127
transform -1 0 5188 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_5
timestamp 1681267127
transform -1 0 4196 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_6
timestamp 1681267127
transform -1 0 3204 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_7
timestamp 1681267127
transform -1 0 2212 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_8
timestamp 1681267127
transform 1 0 7044 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_9
timestamp 1681267127
transform -1 0 1220 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_10
timestamp 1681267127
transform 1 0 6052 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_11
timestamp 1681267127
transform 1 0 5060 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_12
timestamp 1681267127
transform 1 0 1092 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_13
timestamp 1681267127
transform 1 0 2084 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_14
timestamp 1681267127
transform 1 0 3076 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_15
timestamp 1681267127
transform 1 0 4068 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_16
timestamp 1681267127
transform 1 0 9028 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_17
timestamp 1681267127
transform 1 0 10020 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_18
timestamp 1681267127
transform 1 0 11012 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_19
timestamp 1681267127
transform 1 0 12004 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_20
timestamp 1681267127
transform -1 0 9156 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_21
timestamp 1681267127
transform -1 0 10148 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_22
timestamp 1681267127
transform -1 0 11140 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_23
timestamp 1681267127
transform -1 0 12132 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_24
timestamp 1681267127
transform 1 0 12996 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_25
timestamp 1681267127
transform -1 0 13124 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_26
timestamp 1681267127
transform -1 0 13124 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_27
timestamp 1681267127
transform 1 0 12996 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_28
timestamp 1681267127
transform -1 0 12132 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_29
timestamp 1681267127
transform -1 0 11140 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_30
timestamp 1681267127
transform -1 0 10148 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_31
timestamp 1681267127
transform -1 0 9156 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_32
timestamp 1681267127
transform 1 0 12004 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_33
timestamp 1681267127
transform 1 0 11012 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_34
timestamp 1681267127
transform 1 0 10020 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_35
timestamp 1681267127
transform 1 0 9028 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_36
timestamp 1681267127
transform 1 0 4068 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_37
timestamp 1681267127
transform 1 0 3076 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_38
timestamp 1681267127
transform 1 0 2084 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_39
timestamp 1681267127
transform 1 0 1092 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_40
timestamp 1681267127
transform 1 0 5060 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_41
timestamp 1681267127
transform 1 0 6052 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_42
timestamp 1681267127
transform -1 0 1220 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_43
timestamp 1681267127
transform 1 0 7044 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_44
timestamp 1681267127
transform -1 0 2212 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_45
timestamp 1681267127
transform -1 0 3204 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_46
timestamp 1681267127
transform -1 0 4196 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_47
timestamp 1681267127
transform -1 0 5188 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_48
timestamp 1681267127
transform -1 0 6180 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_49
timestamp 1681267127
transform -1 0 7172 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_50
timestamp 1681267127
transform 1 0 8036 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_51
timestamp 1681267127
transform -1 0 8164 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_52
timestamp 1681267127
transform 1 0 734 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_53
timestamp 1681267127
transform -1 0 14401 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_54
timestamp 1681267127
transform 1 0 13988 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_55
timestamp 1681267127
transform 1 0 13988 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_56
timestamp 1681267127
transform -1 0 14401 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_57
timestamp 1681267127
transform 1 0 734 0 1 3152
box 0 0 1 1
use sky130_fd_pr__pfet_01v8__example_55959141808657  sky130_fd_pr__pfet_01v8__example_55959141808657_0
timestamp 1681267127
transform 1 0 14135 0 1 1552
box 0 0 1 1
use sky130_fd_pr__pfet_01v8__example_55959141808657  sky130_fd_pr__pfet_01v8__example_55959141808657_1
timestamp 1681267127
transform 1 0 14135 0 1 3152
box 0 0 1 1
use sky130_fd_pr__pfet_01v8__example_55959141808658  sky130_fd_pr__pfet_01v8__example_55959141808658_0
timestamp 1681267127
transform 1 0 881 0 -1 2552
box 641 0 12546 1
use sky130_fd_pr__pfet_01v8__example_55959141808658  sky130_fd_pr__pfet_01v8__example_55959141808658_1
timestamp 1681267127
transform 1 0 881 0 1 3152
box 641 0 12546 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_0
timestamp 1681267127
transform 1 0 1371 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_1
timestamp 1681267127
transform 1 0 7885 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_2
timestamp 1681267127
transform 1 0 6893 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_3
timestamp 1681267127
transform 1 0 5901 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_4
timestamp 1681267127
transform 1 0 4909 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_5
timestamp 1681267127
transform 1 0 3917 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_6
timestamp 1681267127
transform 1 0 2925 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_7
timestamp 1681267127
transform 1 0 1933 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_8
timestamp 1681267127
transform 1 0 10861 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_9
timestamp 1681267127
transform 1 0 9869 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_10
timestamp 1681267127
transform 1 0 8877 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_11
timestamp 1681267127
transform 1 0 11291 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_12
timestamp 1681267127
transform 1 0 10299 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_13
timestamp 1681267127
transform 1 0 9307 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_14
timestamp 1681267127
transform 1 0 2363 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_15
timestamp 1681267127
transform 1 0 3355 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_16
timestamp 1681267127
transform 1 0 4347 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_17
timestamp 1681267127
transform 1 0 5339 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_18
timestamp 1681267127
transform 1 0 6331 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_19
timestamp 1681267127
transform 1 0 7323 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_20
timestamp 1681267127
transform 1 0 8315 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_21
timestamp 1681267127
transform 1 0 11853 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_22
timestamp 1681267127
transform 1 0 12283 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_23
timestamp 1681267127
transform 1 0 13275 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_24
timestamp 1681267127
transform 1 0 12845 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_25
timestamp 1681267127
transform 1 0 13837 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_26
timestamp 1681267127
transform 1 0 14195 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418085  sky130_fd_pr__via_l1m1_centered__example_559591418085_0
timestamp 1681267127
transform -1 0 14924 0 1 365
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418085  sky130_fd_pr__via_l1m1_centered__example_559591418085_1
timestamp 1681267127
transform -1 0 68 0 1 348
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418086  sky130_fd_pr__via_l1m1_centered__example_559591418086_0
timestamp 1681267127
transform 1 0 941 0 1 1197
box 0 0 1 1
<< properties >>
string GDS_END 5501400
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 4820766
<< end >>
