magic
tech sky130A
magscale 1 2
timestamp 1681267127
<< pwell >>
rect 0 66 756 720
<< nmos >>
rect 194 92 244 694
rect 300 92 350 694
rect 406 92 456 694
rect 512 92 562 694
<< ndiff >>
rect 138 682 194 694
rect 138 648 149 682
rect 183 648 194 682
rect 138 614 194 648
rect 138 580 149 614
rect 183 580 194 614
rect 138 546 194 580
rect 138 512 149 546
rect 183 512 194 546
rect 138 478 194 512
rect 138 444 149 478
rect 183 444 194 478
rect 138 410 194 444
rect 138 376 149 410
rect 183 376 194 410
rect 138 342 194 376
rect 138 308 149 342
rect 183 308 194 342
rect 138 274 194 308
rect 138 240 149 274
rect 183 240 194 274
rect 138 206 194 240
rect 138 172 149 206
rect 183 172 194 206
rect 138 138 194 172
rect 138 104 149 138
rect 183 104 194 138
rect 138 92 194 104
rect 244 682 300 694
rect 244 648 255 682
rect 289 648 300 682
rect 244 614 300 648
rect 244 580 255 614
rect 289 580 300 614
rect 244 546 300 580
rect 244 512 255 546
rect 289 512 300 546
rect 244 478 300 512
rect 244 444 255 478
rect 289 444 300 478
rect 244 410 300 444
rect 244 376 255 410
rect 289 376 300 410
rect 244 342 300 376
rect 244 308 255 342
rect 289 308 300 342
rect 244 274 300 308
rect 244 240 255 274
rect 289 240 300 274
rect 244 206 300 240
rect 244 172 255 206
rect 289 172 300 206
rect 244 138 300 172
rect 244 104 255 138
rect 289 104 300 138
rect 244 92 300 104
rect 350 682 406 694
rect 350 648 361 682
rect 395 648 406 682
rect 350 614 406 648
rect 350 580 361 614
rect 395 580 406 614
rect 350 546 406 580
rect 350 512 361 546
rect 395 512 406 546
rect 350 478 406 512
rect 350 444 361 478
rect 395 444 406 478
rect 350 410 406 444
rect 350 376 361 410
rect 395 376 406 410
rect 350 342 406 376
rect 350 308 361 342
rect 395 308 406 342
rect 350 274 406 308
rect 350 240 361 274
rect 395 240 406 274
rect 350 206 406 240
rect 350 172 361 206
rect 395 172 406 206
rect 350 138 406 172
rect 350 104 361 138
rect 395 104 406 138
rect 350 92 406 104
rect 456 682 512 694
rect 456 648 467 682
rect 501 648 512 682
rect 456 614 512 648
rect 456 580 467 614
rect 501 580 512 614
rect 456 546 512 580
rect 456 512 467 546
rect 501 512 512 546
rect 456 478 512 512
rect 456 444 467 478
rect 501 444 512 478
rect 456 410 512 444
rect 456 376 467 410
rect 501 376 512 410
rect 456 342 512 376
rect 456 308 467 342
rect 501 308 512 342
rect 456 274 512 308
rect 456 240 467 274
rect 501 240 512 274
rect 456 206 512 240
rect 456 172 467 206
rect 501 172 512 206
rect 456 138 512 172
rect 456 104 467 138
rect 501 104 512 138
rect 456 92 512 104
rect 562 682 618 694
rect 562 648 573 682
rect 607 648 618 682
rect 562 614 618 648
rect 562 580 573 614
rect 607 580 618 614
rect 562 546 618 580
rect 562 512 573 546
rect 607 512 618 546
rect 562 478 618 512
rect 562 444 573 478
rect 607 444 618 478
rect 562 410 618 444
rect 562 376 573 410
rect 607 376 618 410
rect 562 342 618 376
rect 562 308 573 342
rect 607 308 618 342
rect 562 274 618 308
rect 562 240 573 274
rect 607 240 618 274
rect 562 206 618 240
rect 562 172 573 206
rect 607 172 618 206
rect 562 138 618 172
rect 562 104 573 138
rect 607 104 618 138
rect 562 92 618 104
<< ndiffc >>
rect 149 648 183 682
rect 149 580 183 614
rect 149 512 183 546
rect 149 444 183 478
rect 149 376 183 410
rect 149 308 183 342
rect 149 240 183 274
rect 149 172 183 206
rect 149 104 183 138
rect 255 648 289 682
rect 255 580 289 614
rect 255 512 289 546
rect 255 444 289 478
rect 255 376 289 410
rect 255 308 289 342
rect 255 240 289 274
rect 255 172 289 206
rect 255 104 289 138
rect 361 648 395 682
rect 361 580 395 614
rect 361 512 395 546
rect 361 444 395 478
rect 361 376 395 410
rect 361 308 395 342
rect 361 240 395 274
rect 361 172 395 206
rect 361 104 395 138
rect 467 648 501 682
rect 467 580 501 614
rect 467 512 501 546
rect 467 444 501 478
rect 467 376 501 410
rect 467 308 501 342
rect 467 240 501 274
rect 467 172 501 206
rect 467 104 501 138
rect 573 648 607 682
rect 573 580 607 614
rect 573 512 607 546
rect 573 444 607 478
rect 573 376 607 410
rect 573 308 607 342
rect 573 240 607 274
rect 573 172 607 206
rect 573 104 607 138
<< psubdiff >>
rect 26 648 84 694
rect 26 614 38 648
rect 72 614 84 648
rect 26 580 84 614
rect 26 546 38 580
rect 72 546 84 580
rect 26 512 84 546
rect 26 478 38 512
rect 72 478 84 512
rect 26 444 84 478
rect 26 410 38 444
rect 72 410 84 444
rect 26 376 84 410
rect 26 342 38 376
rect 72 342 84 376
rect 26 308 84 342
rect 26 274 38 308
rect 72 274 84 308
rect 26 240 84 274
rect 26 206 38 240
rect 72 206 84 240
rect 26 172 84 206
rect 26 138 38 172
rect 72 138 84 172
rect 26 92 84 138
rect 672 648 730 694
rect 672 614 684 648
rect 718 614 730 648
rect 672 580 730 614
rect 672 546 684 580
rect 718 546 730 580
rect 672 512 730 546
rect 672 478 684 512
rect 718 478 730 512
rect 672 444 730 478
rect 672 410 684 444
rect 718 410 730 444
rect 672 376 730 410
rect 672 342 684 376
rect 718 342 730 376
rect 672 308 730 342
rect 672 274 684 308
rect 718 274 730 308
rect 672 240 730 274
rect 672 206 684 240
rect 718 206 730 240
rect 672 172 730 206
rect 672 138 684 172
rect 718 138 730 172
rect 672 92 730 138
<< psubdiffcont >>
rect 38 614 72 648
rect 38 546 72 580
rect 38 478 72 512
rect 38 410 72 444
rect 38 342 72 376
rect 38 274 72 308
rect 38 206 72 240
rect 38 138 72 172
rect 684 614 718 648
rect 684 546 718 580
rect 684 478 718 512
rect 684 410 718 444
rect 684 342 718 376
rect 684 274 718 308
rect 684 206 718 240
rect 684 138 718 172
<< poly >>
rect 175 766 581 786
rect 175 732 191 766
rect 225 732 259 766
rect 293 732 327 766
rect 361 732 395 766
rect 429 732 463 766
rect 497 732 531 766
rect 565 732 581 766
rect 175 716 581 732
rect 175 54 581 70
rect 175 20 191 54
rect 225 20 259 54
rect 293 20 327 54
rect 361 20 395 54
rect 429 20 463 54
rect 497 20 531 54
rect 565 20 581 54
rect 175 0 581 20
<< polycont >>
rect 191 732 225 766
rect 259 732 293 766
rect 327 732 361 766
rect 395 732 429 766
rect 463 732 497 766
rect 531 732 565 766
rect 191 20 225 54
rect 259 20 293 54
rect 327 20 361 54
rect 395 20 429 54
rect 463 20 497 54
rect 531 20 565 54
<< locali >>
rect 175 732 182 766
rect 225 732 254 766
rect 293 732 326 766
rect 361 732 395 766
rect 432 732 463 766
rect 504 732 531 766
rect 576 732 581 766
rect 149 682 183 698
rect 38 662 72 664
rect 38 590 72 614
rect 38 518 72 546
rect 38 446 72 478
rect 38 376 72 410
rect 38 308 72 340
rect 38 240 72 268
rect 38 172 72 196
rect 38 122 72 124
rect 149 614 183 628
rect 149 546 183 556
rect 149 478 183 484
rect 149 410 183 412
rect 149 374 183 376
rect 149 302 183 308
rect 149 230 183 240
rect 149 158 183 172
rect 149 88 183 104
rect 255 682 289 698
rect 255 614 289 628
rect 255 546 289 556
rect 255 478 289 484
rect 255 410 289 412
rect 255 374 289 376
rect 255 302 289 308
rect 255 230 289 240
rect 255 158 289 172
rect 255 88 289 104
rect 361 682 395 698
rect 361 614 395 628
rect 361 546 395 556
rect 361 478 395 484
rect 361 410 395 412
rect 361 374 395 376
rect 361 302 395 308
rect 361 230 395 240
rect 361 158 395 172
rect 361 88 395 104
rect 467 682 501 698
rect 467 614 501 628
rect 467 546 501 556
rect 467 478 501 484
rect 467 410 501 412
rect 467 374 501 376
rect 467 302 501 308
rect 467 230 501 240
rect 467 158 501 172
rect 467 88 501 104
rect 573 682 607 698
rect 573 614 607 628
rect 573 546 607 556
rect 573 478 607 484
rect 573 410 607 412
rect 573 374 607 376
rect 573 302 607 308
rect 573 230 607 240
rect 573 158 607 172
rect 684 662 718 664
rect 684 590 718 614
rect 684 518 718 546
rect 684 446 718 478
rect 684 376 718 410
rect 684 308 718 340
rect 684 240 718 268
rect 684 172 718 196
rect 684 122 718 124
rect 573 88 607 104
rect 175 20 182 54
rect 225 20 254 54
rect 293 20 326 54
rect 361 20 395 54
rect 432 20 463 54
rect 504 20 531 54
rect 576 20 581 54
<< viali >>
rect 182 732 191 766
rect 191 732 216 766
rect 254 732 259 766
rect 259 732 288 766
rect 326 732 327 766
rect 327 732 360 766
rect 398 732 429 766
rect 429 732 432 766
rect 470 732 497 766
rect 497 732 504 766
rect 542 732 565 766
rect 565 732 576 766
rect 38 648 72 662
rect 38 628 72 648
rect 38 580 72 590
rect 38 556 72 580
rect 38 512 72 518
rect 38 484 72 512
rect 38 444 72 446
rect 38 412 72 444
rect 38 342 72 374
rect 38 340 72 342
rect 38 274 72 302
rect 38 268 72 274
rect 38 206 72 230
rect 38 196 72 206
rect 38 138 72 158
rect 38 124 72 138
rect 149 648 183 662
rect 149 628 183 648
rect 149 580 183 590
rect 149 556 183 580
rect 149 512 183 518
rect 149 484 183 512
rect 149 444 183 446
rect 149 412 183 444
rect 149 342 183 374
rect 149 340 183 342
rect 149 274 183 302
rect 149 268 183 274
rect 149 206 183 230
rect 149 196 183 206
rect 149 138 183 158
rect 149 124 183 138
rect 255 648 289 662
rect 255 628 289 648
rect 255 580 289 590
rect 255 556 289 580
rect 255 512 289 518
rect 255 484 289 512
rect 255 444 289 446
rect 255 412 289 444
rect 255 342 289 374
rect 255 340 289 342
rect 255 274 289 302
rect 255 268 289 274
rect 255 206 289 230
rect 255 196 289 206
rect 255 138 289 158
rect 255 124 289 138
rect 361 648 395 662
rect 361 628 395 648
rect 361 580 395 590
rect 361 556 395 580
rect 361 512 395 518
rect 361 484 395 512
rect 361 444 395 446
rect 361 412 395 444
rect 361 342 395 374
rect 361 340 395 342
rect 361 274 395 302
rect 361 268 395 274
rect 361 206 395 230
rect 361 196 395 206
rect 361 138 395 158
rect 361 124 395 138
rect 467 648 501 662
rect 467 628 501 648
rect 467 580 501 590
rect 467 556 501 580
rect 467 512 501 518
rect 467 484 501 512
rect 467 444 501 446
rect 467 412 501 444
rect 467 342 501 374
rect 467 340 501 342
rect 467 274 501 302
rect 467 268 501 274
rect 467 206 501 230
rect 467 196 501 206
rect 467 138 501 158
rect 467 124 501 138
rect 573 648 607 662
rect 573 628 607 648
rect 573 580 607 590
rect 573 556 607 580
rect 573 512 607 518
rect 573 484 607 512
rect 573 444 607 446
rect 573 412 607 444
rect 573 342 607 374
rect 573 340 607 342
rect 573 274 607 302
rect 573 268 607 274
rect 573 206 607 230
rect 573 196 607 206
rect 573 138 607 158
rect 573 124 607 138
rect 684 648 718 662
rect 684 628 718 648
rect 684 580 718 590
rect 684 556 718 580
rect 684 512 718 518
rect 684 484 718 512
rect 684 444 718 446
rect 684 412 718 444
rect 684 342 718 374
rect 684 340 718 342
rect 684 274 718 302
rect 684 268 718 274
rect 684 206 718 230
rect 684 196 718 206
rect 684 138 718 158
rect 684 124 718 138
rect 182 20 191 54
rect 191 20 216 54
rect 254 20 259 54
rect 259 20 288 54
rect 326 20 327 54
rect 327 20 360 54
rect 398 20 429 54
rect 429 20 432 54
rect 470 20 497 54
rect 497 20 504 54
rect 542 20 565 54
rect 565 20 576 54
<< metal1 >>
rect 170 766 588 786
rect 170 732 182 766
rect 216 732 254 766
rect 288 732 326 766
rect 360 732 398 766
rect 432 732 470 766
rect 504 732 542 766
rect 576 732 588 766
rect 170 720 588 732
rect 26 662 84 674
rect 26 628 38 662
rect 72 628 84 662
rect 26 590 84 628
rect 26 556 38 590
rect 72 556 84 590
rect 26 518 84 556
rect 26 484 38 518
rect 72 484 84 518
rect 26 446 84 484
rect 26 412 38 446
rect 72 412 84 446
rect 26 374 84 412
rect 26 340 38 374
rect 72 340 84 374
rect 26 302 84 340
rect 26 268 38 302
rect 72 268 84 302
rect 26 230 84 268
rect 26 196 38 230
rect 72 196 84 230
rect 26 158 84 196
rect 26 124 38 158
rect 72 124 84 158
rect 26 112 84 124
rect 140 662 192 674
rect 140 628 149 662
rect 183 628 192 662
rect 140 590 192 628
rect 140 556 149 590
rect 183 556 192 590
rect 140 518 192 556
rect 140 484 149 518
rect 183 484 192 518
rect 140 446 192 484
rect 140 412 149 446
rect 183 412 192 446
rect 140 374 192 412
rect 140 362 149 374
rect 183 362 192 374
rect 140 302 192 310
rect 140 298 149 302
rect 183 298 192 302
rect 140 234 192 246
rect 140 170 192 182
rect 140 112 192 118
rect 246 668 298 674
rect 246 604 298 616
rect 246 540 298 552
rect 246 484 255 488
rect 289 484 298 488
rect 246 476 298 484
rect 246 412 255 424
rect 289 412 298 424
rect 246 374 298 412
rect 246 340 255 374
rect 289 340 298 374
rect 246 302 298 340
rect 246 268 255 302
rect 289 268 298 302
rect 246 230 298 268
rect 246 196 255 230
rect 289 196 298 230
rect 246 158 298 196
rect 246 124 255 158
rect 289 124 298 158
rect 246 112 298 124
rect 352 662 404 674
rect 352 628 361 662
rect 395 628 404 662
rect 352 590 404 628
rect 352 556 361 590
rect 395 556 404 590
rect 352 518 404 556
rect 352 484 361 518
rect 395 484 404 518
rect 352 446 404 484
rect 352 412 361 446
rect 395 412 404 446
rect 352 374 404 412
rect 352 362 361 374
rect 395 362 404 374
rect 352 302 404 310
rect 352 298 361 302
rect 395 298 404 302
rect 352 234 404 246
rect 352 170 404 182
rect 352 112 404 118
rect 458 668 510 674
rect 458 604 510 616
rect 458 540 510 552
rect 458 484 467 488
rect 501 484 510 488
rect 458 476 510 484
rect 458 412 467 424
rect 501 412 510 424
rect 458 374 510 412
rect 458 340 467 374
rect 501 340 510 374
rect 458 302 510 340
rect 458 268 467 302
rect 501 268 510 302
rect 458 230 510 268
rect 458 196 467 230
rect 501 196 510 230
rect 458 158 510 196
rect 458 124 467 158
rect 501 124 510 158
rect 458 112 510 124
rect 564 662 616 674
rect 564 628 573 662
rect 607 628 616 662
rect 564 590 616 628
rect 564 556 573 590
rect 607 556 616 590
rect 564 518 616 556
rect 564 484 573 518
rect 607 484 616 518
rect 564 446 616 484
rect 564 412 573 446
rect 607 412 616 446
rect 564 374 616 412
rect 564 362 573 374
rect 607 362 616 374
rect 564 302 616 310
rect 564 298 573 302
rect 607 298 616 302
rect 564 234 616 246
rect 564 170 616 182
rect 564 112 616 118
rect 672 662 730 674
rect 672 628 684 662
rect 718 628 730 662
rect 672 590 730 628
rect 672 556 684 590
rect 718 556 730 590
rect 672 518 730 556
rect 672 484 684 518
rect 718 484 730 518
rect 672 446 730 484
rect 672 412 684 446
rect 718 412 730 446
rect 672 374 730 412
rect 672 340 684 374
rect 718 340 730 374
rect 672 302 730 340
rect 672 268 684 302
rect 718 268 730 302
rect 672 230 730 268
rect 672 196 684 230
rect 718 196 730 230
rect 672 158 730 196
rect 672 124 684 158
rect 718 124 730 158
rect 672 112 730 124
rect 170 54 588 66
rect 170 20 182 54
rect 216 20 254 54
rect 288 20 326 54
rect 360 20 398 54
rect 432 20 470 54
rect 504 20 542 54
rect 576 20 588 54
rect 170 0 588 20
<< via1 >>
rect 140 340 149 362
rect 149 340 183 362
rect 183 340 192 362
rect 140 310 192 340
rect 140 268 149 298
rect 149 268 183 298
rect 183 268 192 298
rect 140 246 192 268
rect 140 230 192 234
rect 140 196 149 230
rect 149 196 183 230
rect 183 196 192 230
rect 140 182 192 196
rect 140 158 192 170
rect 140 124 149 158
rect 149 124 183 158
rect 183 124 192 158
rect 140 118 192 124
rect 246 662 298 668
rect 246 628 255 662
rect 255 628 289 662
rect 289 628 298 662
rect 246 616 298 628
rect 246 590 298 604
rect 246 556 255 590
rect 255 556 289 590
rect 289 556 298 590
rect 246 552 298 556
rect 246 518 298 540
rect 246 488 255 518
rect 255 488 289 518
rect 289 488 298 518
rect 246 446 298 476
rect 246 424 255 446
rect 255 424 289 446
rect 289 424 298 446
rect 352 340 361 362
rect 361 340 395 362
rect 395 340 404 362
rect 352 310 404 340
rect 352 268 361 298
rect 361 268 395 298
rect 395 268 404 298
rect 352 246 404 268
rect 352 230 404 234
rect 352 196 361 230
rect 361 196 395 230
rect 395 196 404 230
rect 352 182 404 196
rect 352 158 404 170
rect 352 124 361 158
rect 361 124 395 158
rect 395 124 404 158
rect 352 118 404 124
rect 458 662 510 668
rect 458 628 467 662
rect 467 628 501 662
rect 501 628 510 662
rect 458 616 510 628
rect 458 590 510 604
rect 458 556 467 590
rect 467 556 501 590
rect 501 556 510 590
rect 458 552 510 556
rect 458 518 510 540
rect 458 488 467 518
rect 467 488 501 518
rect 501 488 510 518
rect 458 446 510 476
rect 458 424 467 446
rect 467 424 501 446
rect 501 424 510 446
rect 564 340 573 362
rect 573 340 607 362
rect 607 340 616 362
rect 564 310 616 340
rect 564 268 573 298
rect 573 268 607 298
rect 607 268 616 298
rect 564 246 616 268
rect 564 230 616 234
rect 564 196 573 230
rect 573 196 607 230
rect 607 196 616 230
rect 564 182 616 196
rect 564 158 616 170
rect 564 124 573 158
rect 573 124 607 158
rect 607 124 616 158
rect 564 118 616 124
<< metal2 >>
rect 0 668 756 674
rect 0 616 246 668
rect 298 616 458 668
rect 510 616 756 668
rect 0 604 756 616
rect 0 552 246 604
rect 298 552 458 604
rect 510 552 756 604
rect 0 540 756 552
rect 0 488 246 540
rect 298 488 458 540
rect 510 488 756 540
rect 0 476 756 488
rect 0 424 246 476
rect 298 424 458 476
rect 510 424 756 476
rect 0 418 756 424
rect 0 362 756 368
rect 0 310 140 362
rect 192 310 352 362
rect 404 310 564 362
rect 616 310 756 362
rect 0 298 756 310
rect 0 246 140 298
rect 192 246 352 298
rect 404 246 564 298
rect 616 246 756 298
rect 0 234 756 246
rect 0 182 140 234
rect 192 182 352 234
rect 404 182 564 234
rect 616 182 756 234
rect 0 170 756 182
rect 0 118 140 170
rect 192 118 352 170
rect 404 118 564 170
rect 616 118 756 170
rect 0 112 756 118
<< labels >>
flabel comment s 166 393 166 393 0 FreeSans 300 0 0 0 S
flabel comment s 272 393 272 393 0 FreeSans 300 0 0 0 S
flabel comment s 378 393 378 393 0 FreeSans 300 0 0 0 S
flabel comment s 484 393 484 393 0 FreeSans 300 0 0 0 S
flabel comment s 166 393 166 393 0 FreeSans 300 0 0 0 S
flabel comment s 272 393 272 393 0 FreeSans 300 0 0 0 D
flabel comment s 378 393 378 393 0 FreeSans 300 0 0 0 S
flabel comment s 484 393 484 393 0 FreeSans 300 0 0 0 D
flabel comment s 590 393 590 393 0 FreeSans 300 0 0 0 S
flabel metal2 s 3 491 22 561 0 FreeSans 400 90 0 0 DRAIN
port 2 nsew
flabel metal2 s 3 180 24 244 0 FreeSans 400 90 0 0 SOURCE
port 3 nsew
flabel metal1 s 288 24 370 49 0 FreeSans 400 0 0 0 GATE
port 4 nsew
flabel metal1 s 347 737 429 762 0 FreeSans 400 0 0 0 GATE
port 4 nsew
flabel metal1 s 51 544 51 544 7 FreeSans 400 90 0 0 SUBSTRATE
flabel metal1 s 700 523 700 523 7 FreeSans 400 90 0 0 SUBSTRATE
<< properties >>
string GDS_END 5073924
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 5058106
<< end >>
