magic
tech sky130A
magscale 1 2
timestamp 1681267127
use sky130_fd_pr__hvdfl1sd2__example_55959141808143  sky130_fd_pr__hvdfl1sd2__example_55959141808143_0
timestamp 1681267127
transform 1 0 100 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808143  sky130_fd_pr__hvdfl1sd2__example_55959141808143_1
timestamp 1681267127
transform 1 0 256 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808102  sky130_fd_pr__hvdfl1sd__example_55959141808102_0
timestamp 1681267127
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808102  sky130_fd_pr__hvdfl1sd__example_55959141808102_1
timestamp 1681267127
transform 1 0 412 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 7310790
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 7308700
<< end >>
