magic
tech sky130A
magscale 1 2
timestamp 1681267127
<< nwell >>
rect 2774 4256 3850 4424
rect 3682 3218 3850 4256
rect 2774 3050 3850 3218
<< pwell >>
rect 3048 3278 3622 4196
<< mvnmos >>
rect 3235 3462 3435 4062
<< mvndiff >>
rect 3182 4050 3235 4062
rect 3182 4016 3190 4050
rect 3224 4016 3235 4050
rect 3182 3982 3235 4016
rect 3182 3948 3190 3982
rect 3224 3948 3235 3982
rect 3182 3914 3235 3948
rect 3182 3880 3190 3914
rect 3224 3880 3235 3914
rect 3182 3846 3235 3880
rect 3182 3812 3190 3846
rect 3224 3812 3235 3846
rect 3182 3778 3235 3812
rect 3182 3744 3190 3778
rect 3224 3744 3235 3778
rect 3182 3710 3235 3744
rect 3182 3676 3190 3710
rect 3224 3676 3235 3710
rect 3182 3642 3235 3676
rect 3182 3608 3190 3642
rect 3224 3608 3235 3642
rect 3182 3574 3235 3608
rect 3182 3540 3190 3574
rect 3224 3540 3235 3574
rect 3182 3462 3235 3540
rect 3435 4050 3488 4062
rect 3435 4016 3446 4050
rect 3480 4016 3488 4050
rect 3435 3982 3488 4016
rect 3435 3948 3446 3982
rect 3480 3948 3488 3982
rect 3435 3914 3488 3948
rect 3435 3880 3446 3914
rect 3480 3880 3488 3914
rect 3435 3846 3488 3880
rect 3435 3812 3446 3846
rect 3480 3812 3488 3846
rect 3435 3778 3488 3812
rect 3435 3744 3446 3778
rect 3480 3744 3488 3778
rect 3435 3710 3488 3744
rect 3435 3676 3446 3710
rect 3480 3676 3488 3710
rect 3435 3642 3488 3676
rect 3435 3608 3446 3642
rect 3480 3608 3488 3642
rect 3435 3574 3488 3608
rect 3435 3540 3446 3574
rect 3480 3540 3488 3574
rect 3435 3462 3488 3540
<< mvndiffc >>
rect 3190 4016 3224 4050
rect 3190 3948 3224 3982
rect 3190 3880 3224 3914
rect 3190 3812 3224 3846
rect 3190 3744 3224 3778
rect 3190 3676 3224 3710
rect 3190 3608 3224 3642
rect 3190 3540 3224 3574
rect 3446 4016 3480 4050
rect 3446 3948 3480 3982
rect 3446 3880 3480 3914
rect 3446 3812 3480 3846
rect 3446 3744 3480 3778
rect 3446 3676 3480 3710
rect 3446 3608 3480 3642
rect 3446 3540 3480 3574
<< mvpsubdiff >>
rect 3074 4136 3188 4170
rect 3222 4136 3256 4170
rect 3290 4136 3324 4170
rect 3358 4136 3392 4170
rect 3426 4136 3460 4170
rect 3494 4136 3528 4170
rect 3074 4068 3108 4102
rect 3562 4068 3596 4170
rect 3074 4000 3108 4034
rect 3074 3932 3108 3966
rect 3074 3864 3108 3898
rect 3074 3796 3108 3830
rect 3074 3728 3108 3762
rect 3074 3660 3108 3694
rect 3074 3592 3108 3626
rect 3074 3524 3108 3558
rect 3074 3456 3108 3490
rect 3562 4000 3596 4034
rect 3562 3932 3596 3966
rect 3562 3864 3596 3898
rect 3562 3796 3596 3830
rect 3562 3728 3596 3762
rect 3562 3660 3596 3694
rect 3562 3592 3596 3626
rect 3562 3524 3596 3558
rect 3074 3304 3108 3422
rect 3562 3372 3596 3490
rect 3142 3304 3176 3338
rect 3210 3304 3244 3338
rect 3278 3304 3312 3338
rect 3346 3304 3380 3338
rect 3414 3304 3448 3338
rect 3482 3304 3596 3338
<< mvnsubdiff >>
rect 2917 4322 2941 4356
rect 2975 4322 3012 4356
rect 3046 4322 3083 4356
rect 3117 4322 3154 4356
rect 3188 4322 3225 4356
rect 3259 4322 3296 4356
rect 3330 4322 3367 4356
rect 3401 4322 3438 4356
rect 3472 4322 3509 4356
rect 3543 4322 3580 4356
rect 3614 4322 3652 4356
rect 3686 4322 3724 4356
rect 3758 4322 3782 4356
rect 3748 4264 3782 4322
rect 3748 4196 3782 4230
rect 3748 4128 3782 4162
rect 3748 4060 3782 4094
rect 3748 3992 3782 4026
rect 3748 3924 3782 3958
rect 3748 3856 3782 3890
rect 3748 3788 3782 3822
rect 3748 3720 3782 3754
rect 3748 3652 3782 3686
rect 3748 3584 3782 3618
rect 3748 3516 3782 3550
rect 3748 3448 3782 3482
rect 3748 3380 3782 3414
rect 3748 3312 3782 3346
rect 3748 3244 3782 3278
rect 3748 3176 3782 3210
rect 2919 3118 2943 3152
rect 2977 3118 3014 3152
rect 3048 3118 3085 3152
rect 3119 3118 3156 3152
rect 3190 3118 3227 3152
rect 3261 3118 3298 3152
rect 3332 3118 3369 3152
rect 3403 3118 3440 3152
rect 3474 3118 3511 3152
rect 3545 3118 3582 3152
rect 3616 3118 3652 3152
rect 3686 3142 3748 3152
rect 3686 3118 3782 3142
<< mvpsubdiffcont >>
rect 3188 4136 3222 4170
rect 3256 4136 3290 4170
rect 3324 4136 3358 4170
rect 3392 4136 3426 4170
rect 3460 4136 3494 4170
rect 3528 4136 3562 4170
rect 3074 4102 3108 4136
rect 3074 4034 3108 4068
rect 3074 3966 3108 4000
rect 3074 3898 3108 3932
rect 3074 3830 3108 3864
rect 3074 3762 3108 3796
rect 3074 3694 3108 3728
rect 3074 3626 3108 3660
rect 3074 3558 3108 3592
rect 3074 3490 3108 3524
rect 3562 4034 3596 4068
rect 3562 3966 3596 4000
rect 3562 3898 3596 3932
rect 3562 3830 3596 3864
rect 3562 3762 3596 3796
rect 3562 3694 3596 3728
rect 3562 3626 3596 3660
rect 3562 3558 3596 3592
rect 3562 3490 3596 3524
rect 3074 3422 3108 3456
rect 3562 3338 3596 3372
rect 3108 3304 3142 3338
rect 3176 3304 3210 3338
rect 3244 3304 3278 3338
rect 3312 3304 3346 3338
rect 3380 3304 3414 3338
rect 3448 3304 3482 3338
<< mvnsubdiffcont >>
rect 2941 4322 2975 4356
rect 3012 4322 3046 4356
rect 3083 4322 3117 4356
rect 3154 4322 3188 4356
rect 3225 4322 3259 4356
rect 3296 4322 3330 4356
rect 3367 4322 3401 4356
rect 3438 4322 3472 4356
rect 3509 4322 3543 4356
rect 3580 4322 3614 4356
rect 3652 4322 3686 4356
rect 3724 4322 3758 4356
rect 3748 4230 3782 4264
rect 3748 4162 3782 4196
rect 3748 4094 3782 4128
rect 3748 4026 3782 4060
rect 3748 3958 3782 3992
rect 3748 3890 3782 3924
rect 3748 3822 3782 3856
rect 3748 3754 3782 3788
rect 3748 3686 3782 3720
rect 3748 3618 3782 3652
rect 3748 3550 3782 3584
rect 3748 3482 3782 3516
rect 3748 3414 3782 3448
rect 3748 3346 3782 3380
rect 3748 3278 3782 3312
rect 3748 3210 3782 3244
rect 2943 3118 2977 3152
rect 3014 3118 3048 3152
rect 3085 3118 3119 3152
rect 3156 3118 3190 3152
rect 3227 3118 3261 3152
rect 3298 3118 3332 3152
rect 3369 3118 3403 3152
rect 3440 3118 3474 3152
rect 3511 3118 3545 3152
rect 3582 3118 3616 3152
rect 3652 3118 3686 3152
rect 3748 3142 3782 3176
<< poly >>
rect 3235 3436 3435 3462
rect 3235 3420 3437 3436
rect 3235 3386 3251 3420
rect 3285 3386 3319 3420
rect 3353 3386 3387 3420
rect 3421 3386 3437 3420
rect 3235 3370 3437 3386
<< polycont >>
rect 3251 3386 3285 3420
rect 3319 3386 3353 3420
rect 3387 3386 3421 3420
<< locali >>
rect 2272 4572 2310 4606
rect 2344 4572 2382 4606
rect 2917 4322 2941 4356
rect 3009 4322 3012 4356
rect 3046 4322 3047 4356
rect 3081 4322 3083 4356
rect 3117 4322 3119 4356
rect 3153 4322 3154 4356
rect 3188 4322 3191 4356
rect 3259 4322 3263 4356
rect 3330 4322 3335 4356
rect 3401 4322 3407 4356
rect 3472 4322 3479 4356
rect 3543 4322 3551 4356
rect 3614 4322 3623 4356
rect 3686 4322 3695 4356
rect 3758 4322 3782 4356
rect 3748 4264 3782 4322
rect 3748 4196 3782 4211
rect 3074 4152 3169 4170
rect 3108 4136 3169 4152
rect 3222 4136 3241 4170
rect 3290 4136 3313 4170
rect 3358 4136 3385 4170
rect 3426 4136 3457 4170
rect 3494 4136 3528 4170
rect 3074 4080 3108 4102
rect 3562 4098 3596 4136
rect 3074 4008 3108 4034
rect 3074 3936 3108 3966
rect 3074 3864 3108 3898
rect 3074 3796 3108 3830
rect 3074 3728 3108 3758
rect 3074 3660 3108 3686
rect 3074 3592 3108 3614
rect 3074 3524 3108 3542
rect 3190 4063 3224 4066
rect 3190 3991 3224 4016
rect 3190 3919 3224 3948
rect 3190 3847 3224 3880
rect 3190 3778 3224 3812
rect 3190 3710 3224 3741
rect 3190 3642 3224 3669
rect 3190 3574 3224 3597
rect 3190 3524 3224 3525
rect 3446 4004 3480 4016
rect 3446 3914 3480 3948
rect 3446 3846 3480 3880
rect 3446 3797 3480 3812
rect 3446 3725 3480 3744
rect 3446 3653 3480 3676
rect 3446 3581 3480 3608
rect 3446 3524 3480 3540
rect 3562 4026 3596 4034
rect 3562 3932 3596 3966
rect 3562 3864 3596 3898
rect 3562 3796 3596 3804
rect 3562 3728 3596 3732
rect 3562 3592 3596 3626
rect 3562 3524 3596 3558
rect 3074 3456 3108 3470
rect 3562 3448 3596 3486
rect 3074 3360 3108 3398
rect 3235 3386 3251 3420
rect 3317 3386 3319 3420
rect 3353 3386 3355 3420
rect 3421 3386 3437 3420
rect 3562 3376 3596 3414
rect 3074 3304 3108 3326
rect 3142 3304 3164 3338
rect 3210 3304 3244 3338
rect 3280 3304 3312 3338
rect 3362 3304 3380 3338
rect 3443 3304 3448 3338
rect 3482 3304 3490 3338
rect 3524 3304 3596 3338
rect 3748 4128 3782 4139
rect 3748 4060 3782 4067
rect 3748 3992 3782 3995
rect 3748 3924 3782 3958
rect 3748 3856 3782 3890
rect 3748 3788 3782 3804
rect 3748 3720 3782 3732
rect 3748 3652 3782 3660
rect 3748 3584 3782 3618
rect 3748 3516 3782 3550
rect 3748 3448 3782 3474
rect 3748 3380 3782 3402
rect 3748 3312 3782 3330
rect 3748 3244 3782 3258
rect 3748 3176 3782 3186
rect 2919 3118 2943 3152
rect 3006 3118 3014 3152
rect 3078 3118 3085 3152
rect 3150 3118 3156 3152
rect 3222 3118 3227 3152
rect 3294 3118 3298 3152
rect 3366 3118 3369 3152
rect 3403 3118 3404 3152
rect 3438 3118 3440 3152
rect 3474 3118 3476 3152
rect 3510 3118 3511 3152
rect 3545 3118 3548 3152
rect 3616 3118 3620 3152
rect 3686 3118 3692 3152
rect 3726 3142 3748 3152
rect 3726 3118 3782 3142
rect 2272 246 2310 280
rect 2344 246 2382 280
<< viali >>
rect 2238 4572 2272 4606
rect 2310 4572 2344 4606
rect 2382 4572 2416 4606
rect 2975 4322 3009 4356
rect 3047 4322 3081 4356
rect 3119 4322 3153 4356
rect 3191 4322 3225 4356
rect 3263 4322 3296 4356
rect 3296 4322 3297 4356
rect 3335 4322 3367 4356
rect 3367 4322 3369 4356
rect 3407 4322 3438 4356
rect 3438 4322 3441 4356
rect 3479 4322 3509 4356
rect 3509 4322 3513 4356
rect 3551 4322 3580 4356
rect 3580 4322 3585 4356
rect 3623 4322 3652 4356
rect 3652 4322 3657 4356
rect 3695 4322 3724 4356
rect 3724 4322 3729 4356
rect 3748 4230 3782 4245
rect 3748 4211 3782 4230
rect 3074 4136 3108 4152
rect 3169 4136 3188 4170
rect 3188 4136 3203 4170
rect 3241 4136 3256 4170
rect 3256 4136 3275 4170
rect 3313 4136 3324 4170
rect 3324 4136 3347 4170
rect 3385 4136 3392 4170
rect 3392 4136 3419 4170
rect 3457 4136 3460 4170
rect 3460 4136 3491 4170
rect 3562 4136 3596 4170
rect 3074 4118 3108 4136
rect 3074 4068 3108 4080
rect 3074 4046 3108 4068
rect 3074 4000 3108 4008
rect 3074 3974 3108 4000
rect 3074 3932 3108 3936
rect 3074 3902 3108 3932
rect 3074 3830 3108 3864
rect 3074 3762 3108 3792
rect 3074 3758 3108 3762
rect 3074 3694 3108 3720
rect 3074 3686 3108 3694
rect 3074 3626 3108 3648
rect 3074 3614 3108 3626
rect 3074 3558 3108 3576
rect 3074 3542 3108 3558
rect 3190 4050 3224 4063
rect 3190 4029 3224 4050
rect 3190 3982 3224 3991
rect 3190 3957 3224 3982
rect 3190 3914 3224 3919
rect 3190 3885 3224 3914
rect 3190 3846 3224 3847
rect 3190 3813 3224 3846
rect 3190 3744 3224 3775
rect 3190 3741 3224 3744
rect 3190 3676 3224 3703
rect 3190 3669 3224 3676
rect 3190 3608 3224 3631
rect 3190 3597 3224 3608
rect 3190 3540 3224 3559
rect 3190 3525 3224 3540
rect 3446 4050 3480 4076
rect 3446 4042 3480 4050
rect 3446 3982 3480 4004
rect 3446 3970 3480 3982
rect 3446 3778 3480 3797
rect 3446 3763 3480 3778
rect 3446 3710 3480 3725
rect 3446 3691 3480 3710
rect 3446 3642 3480 3653
rect 3446 3619 3480 3642
rect 3446 3574 3480 3581
rect 3446 3547 3480 3574
rect 3562 4068 3596 4098
rect 3562 4064 3596 4068
rect 3562 4000 3596 4026
rect 3562 3992 3596 4000
rect 3562 3830 3596 3838
rect 3562 3804 3596 3830
rect 3562 3762 3596 3766
rect 3562 3732 3596 3762
rect 3562 3660 3596 3694
rect 3074 3490 3108 3504
rect 3074 3470 3108 3490
rect 3074 3422 3108 3432
rect 3074 3398 3108 3422
rect 3562 3490 3596 3520
rect 3562 3486 3596 3490
rect 3283 3386 3285 3420
rect 3285 3386 3317 3420
rect 3355 3386 3387 3420
rect 3387 3386 3389 3420
rect 3562 3414 3596 3448
rect 3074 3326 3108 3360
rect 3562 3372 3596 3376
rect 3562 3342 3596 3372
rect 3164 3304 3176 3338
rect 3176 3304 3198 3338
rect 3246 3304 3278 3338
rect 3278 3304 3280 3338
rect 3328 3304 3346 3338
rect 3346 3304 3362 3338
rect 3409 3304 3414 3338
rect 3414 3304 3443 3338
rect 3490 3304 3524 3338
rect 3748 4162 3782 4173
rect 3748 4139 3782 4162
rect 3748 4094 3782 4101
rect 3748 4067 3782 4094
rect 3748 4026 3782 4029
rect 3748 3995 3782 4026
rect 3748 3822 3782 3838
rect 3748 3804 3782 3822
rect 3748 3754 3782 3766
rect 3748 3732 3782 3754
rect 3748 3686 3782 3694
rect 3748 3660 3782 3686
rect 3748 3482 3782 3508
rect 3748 3474 3782 3482
rect 3748 3414 3782 3436
rect 3748 3402 3782 3414
rect 3748 3346 3782 3364
rect 3748 3330 3782 3346
rect 3748 3278 3782 3292
rect 3748 3258 3782 3278
rect 3748 3210 3782 3220
rect 3748 3186 3782 3210
rect 2972 3118 2977 3152
rect 2977 3118 3006 3152
rect 3044 3118 3048 3152
rect 3048 3118 3078 3152
rect 3116 3118 3119 3152
rect 3119 3118 3150 3152
rect 3188 3118 3190 3152
rect 3190 3118 3222 3152
rect 3260 3118 3261 3152
rect 3261 3118 3294 3152
rect 3332 3118 3366 3152
rect 3404 3118 3438 3152
rect 3476 3118 3510 3152
rect 3548 3118 3582 3152
rect 3620 3118 3652 3152
rect 3652 3118 3654 3152
rect 3692 3118 3726 3152
rect 2238 246 2272 280
rect 2310 246 2344 280
rect 2382 246 2416 280
<< metal1 >>
rect 2455 4626 4014 4651
rect 276 4510 282 4626
rect 590 4510 596 4626
rect 1468 4510 1474 4626
rect 1590 4510 1596 4626
rect 2230 4510 2236 4626
rect 2416 4510 2422 4626
rect 2455 4510 2461 4626
rect 2705 4510 4014 4626
rect 2455 4508 4014 4510
rect 2776 4449 4014 4508
rect 2902 4365 4014 4449
rect 2902 4356 3794 4365
rect 2902 4348 2975 4356
rect 2920 4322 2975 4348
rect 3009 4322 3047 4356
rect 3081 4322 3119 4356
rect 3153 4322 3191 4356
rect 3225 4322 3263 4356
rect 3297 4322 3335 4356
rect 3369 4322 3407 4356
rect 3441 4322 3479 4356
rect 3513 4322 3551 4356
rect 3585 4322 3623 4356
rect 3657 4322 3695 4356
rect 3729 4322 3794 4356
rect 2920 4316 3794 4322
tri 2920 4278 2958 4316 nw
tri 3678 4278 3716 4316 ne
rect 3716 4245 3794 4316
tri 3794 4306 3853 4365 nw
rect 3716 4211 3748 4245
rect 3782 4211 3794 4245
rect 440 4066 446 4182
rect 562 4066 568 4182
rect 1158 4066 1164 4182
rect 1280 4066 1286 4182
rect 1780 4066 1786 4182
rect 1902 4066 1908 4182
rect 2495 4066 2501 4182
rect 2617 4066 2623 4182
rect 2948 4066 2959 4182
rect 3075 4170 3608 4182
rect 3075 4152 3169 4170
rect 3108 4136 3169 4152
rect 3203 4136 3241 4170
rect 3275 4136 3313 4170
rect 3347 4136 3385 4170
rect 3419 4136 3457 4170
rect 3491 4136 3562 4170
rect 3596 4136 3608 4170
rect 3108 4130 3608 4136
rect 3108 4118 3123 4130
rect 3075 4101 3123 4118
tri 3123 4101 3152 4130 nw
tri 3518 4101 3547 4130 ne
rect 3547 4101 3608 4130
rect 3075 4098 3120 4101
tri 3120 4098 3123 4101 nw
tri 3547 4098 3550 4101 ne
rect 3550 4098 3608 4101
rect 3075 4080 3114 4098
tri 3114 4092 3120 4098 nw
tri 3550 4092 3556 4098 ne
rect 2948 4046 3074 4066
rect 3108 4046 3114 4080
rect 3437 4080 3489 4088
rect 645 4032 825 4038
rect 645 3910 825 3916
rect 1977 4032 2157 4038
rect 1977 3910 2157 3916
rect 2948 4008 3114 4046
rect 2948 3974 3074 4008
rect 3108 3974 3114 4008
rect 2948 3936 3114 3974
rect 2948 3902 3074 3936
rect 3108 3902 3114 3936
rect 440 3766 446 3882
rect 562 3766 568 3882
rect 1159 3766 1165 3882
rect 1281 3766 1287 3882
rect 1775 3766 1781 3882
rect 1897 3766 1903 3882
rect 2495 3766 2501 3882
rect 2617 3766 2623 3882
rect 2948 3875 3114 3902
rect 899 3005 905 3616
tri 838 2923 895 2980 se
rect 895 2924 905 3005
rect 1085 3005 1091 3616
rect 1131 3610 1309 3616
rect 1131 3110 1162 3610
rect 1278 3110 1309 3610
rect 1131 3097 1309 3110
rect 1131 3045 1162 3097
rect 1214 3045 1226 3097
rect 1278 3045 1309 3097
rect 1131 3032 1309 3045
rect 1085 2950 1095 3005
rect 1085 2924 1091 2950
tri 1091 2946 1095 2950 nw
rect 1131 2980 1162 3032
rect 1214 2980 1226 3032
rect 1278 2980 1309 3032
rect 1131 2967 1309 2980
rect 895 2923 1068 2924
tri 1068 2923 1069 2924 nw
rect 895 2892 1021 2923
rect 197 2403 223 2452
rect 826 1944 832 2892
rect 948 2876 1021 2892
tri 1021 2876 1068 2923 nw
rect 1131 2915 1162 2967
rect 1214 2915 1226 2967
rect 1278 2915 1309 2967
rect 1131 2902 1309 2915
rect 948 1976 954 2876
tri 964 2819 1021 2876 nw
rect 1131 2850 1162 2902
rect 1214 2850 1226 2902
rect 1278 2850 1309 2902
rect 1131 2837 1309 2850
rect 1131 2785 1162 2837
rect 1214 2785 1226 2837
rect 1278 2785 1309 2837
rect 1131 2772 1309 2785
rect 1131 2720 1162 2772
rect 1214 2720 1226 2772
rect 1278 2720 1309 2772
rect 1131 2714 1309 2720
rect 1753 3610 1931 3616
rect 1753 3110 1784 3610
rect 1900 3110 1931 3610
rect 2948 3247 2954 3875
rect 3070 3864 3114 3875
rect 3070 3830 3074 3864
rect 3108 3830 3114 3864
rect 3070 3792 3114 3830
rect 3070 3758 3074 3792
rect 3108 3758 3114 3792
rect 3070 3720 3114 3758
rect 3070 3686 3074 3720
rect 3108 3686 3114 3720
rect 3070 3648 3114 3686
rect 3070 3614 3074 3648
rect 3108 3614 3114 3648
rect 3070 3576 3114 3614
rect 3070 3542 3074 3576
rect 3108 3542 3114 3576
rect 3070 3504 3114 3542
rect 3181 4072 3233 4078
rect 3181 4008 3233 4020
rect 3437 4016 3489 4028
rect 3437 3958 3489 3964
rect 3556 4080 3562 4098
rect 3596 4080 3608 4098
rect 3556 4026 3608 4028
rect 3556 4016 3562 4026
rect 3596 4016 3608 4026
rect 3556 3958 3608 3964
rect 3716 4173 3794 4211
rect 3716 4153 3748 4173
rect 3782 4139 3794 4173
rect 3768 4101 3794 4139
rect 3716 4089 3748 4101
rect 3782 4088 3794 4101
tri 3794 4088 3832 4126 sw
rect 3782 4067 4014 4088
rect 3768 4037 4014 4067
rect 3716 4029 4014 4037
rect 3716 4025 3748 4029
rect 3782 3995 4014 4029
rect 3768 3973 4014 3995
rect 3716 3958 4014 3973
rect 3181 3944 3233 3956
tri 3233 3930 3258 3955 sw
rect 3233 3892 4014 3930
rect 3181 3885 3190 3892
rect 3224 3885 4014 3892
rect 3181 3880 4014 3885
rect 3233 3878 4014 3880
tri 3233 3853 3258 3878 nw
rect 3181 3816 3190 3828
rect 3224 3816 3233 3828
rect 3556 3838 3608 3850
rect 3181 3752 3190 3764
rect 3224 3752 3233 3764
rect 3181 3669 3190 3700
rect 3224 3669 3233 3700
rect 3181 3631 3233 3669
rect 3181 3597 3190 3631
rect 3224 3597 3233 3631
rect 3181 3559 3233 3597
rect 3181 3525 3190 3559
rect 3224 3525 3233 3559
rect 3181 3513 3233 3525
rect 3437 3811 3489 3817
rect 3437 3747 3489 3759
rect 3437 3691 3446 3695
rect 3480 3691 3489 3695
rect 3437 3683 3489 3691
rect 3556 3774 3608 3786
rect 3556 3710 3608 3722
rect 3556 3648 3608 3658
rect 3716 3839 3794 3850
rect 3768 3838 3794 3839
rect 3782 3804 3794 3838
rect 3768 3787 3794 3804
rect 3716 3775 3794 3787
rect 3768 3766 3794 3775
rect 3782 3732 3794 3766
rect 3768 3723 3794 3732
rect 3716 3711 3794 3723
rect 3768 3694 3794 3711
rect 3782 3660 3794 3694
rect 3768 3659 3794 3660
rect 3716 3648 3794 3659
rect 3437 3619 3446 3631
rect 3480 3620 3489 3631
tri 3489 3620 3514 3645 sw
rect 3480 3619 4014 3620
rect 3489 3568 4014 3619
rect 3437 3555 3446 3567
rect 3480 3555 3489 3567
rect 3070 3470 3074 3504
rect 3108 3470 3114 3504
tri 3489 3543 3514 3568 nw
rect 3437 3497 3489 3503
rect 3556 3533 3608 3540
rect 3070 3432 3114 3470
rect 3070 3398 3074 3432
rect 3108 3398 3114 3432
rect 3556 3469 3608 3481
rect 3070 3377 3114 3398
tri 3114 3377 3119 3382 sw
rect 3271 3377 3278 3429
rect 3330 3377 3342 3429
rect 3394 3377 3401 3429
rect 3556 3414 3562 3417
rect 3596 3414 3608 3417
rect 3556 3405 3608 3414
tri 3551 3377 3556 3382 se
rect 3070 3376 3119 3377
tri 3119 3376 3120 3377 sw
tri 3550 3376 3551 3377 se
rect 3551 3376 3556 3377
rect 3070 3360 3120 3376
rect 3070 3326 3074 3360
rect 3108 3344 3120 3360
tri 3120 3344 3152 3376 sw
tri 3518 3344 3550 3376 se
rect 3550 3353 3556 3376
rect 3550 3344 3562 3353
rect 3108 3342 3562 3344
rect 3596 3342 3608 3353
rect 3108 3338 3608 3342
rect 3108 3326 3164 3338
rect 3070 3304 3164 3326
rect 3198 3304 3246 3338
rect 3280 3304 3328 3338
rect 3362 3304 3409 3338
rect 3443 3304 3490 3338
rect 3524 3304 3608 3338
rect 3070 3298 3608 3304
rect 3716 3527 3794 3533
rect 3768 3508 3794 3527
rect 3716 3474 3748 3475
rect 3782 3474 3794 3508
rect 3716 3463 3794 3474
rect 3768 3436 3794 3463
rect 3716 3402 3748 3411
rect 3782 3402 3794 3436
rect 3716 3399 3794 3402
rect 3768 3392 3794 3399
tri 3794 3392 3832 3430 sw
rect 3768 3364 4014 3392
rect 3716 3335 3748 3347
rect 3782 3330 4014 3364
rect 3070 3292 3108 3298
tri 3108 3292 3114 3298 nw
rect 3768 3292 4014 3330
rect 3070 3247 3076 3292
tri 3076 3260 3108 3292 nw
rect 3716 3271 3748 3283
rect 2948 3241 3076 3247
rect 3782 3264 4014 3292
rect 3782 3260 3828 3264
tri 3828 3260 3832 3264 nw
rect 3782 3258 3820 3260
rect 3768 3252 3820 3258
tri 3820 3252 3828 3260 nw
rect 3768 3220 3794 3252
tri 3794 3226 3820 3252 nw
rect 3716 3207 3748 3219
tri 3706 3186 3716 3196 se
rect 3782 3186 3794 3220
tri 3703 3183 3706 3186 se
rect 3706 3183 3716 3186
rect 1753 3097 1931 3110
rect 1753 3045 1784 3097
rect 1836 3045 1848 3097
rect 1900 3045 1931 3097
tri 2920 3158 2945 3183 sw
tri 3678 3158 3703 3183 se
rect 3703 3158 3716 3183
rect 2920 3155 3716 3158
rect 3768 3155 3794 3186
rect 2920 3152 3794 3155
rect 2920 3118 2972 3152
rect 3006 3118 3044 3152
rect 3078 3118 3116 3152
rect 3150 3118 3188 3152
rect 3222 3118 3260 3152
rect 3294 3118 3332 3152
rect 3366 3118 3404 3152
rect 3438 3118 3476 3152
rect 3510 3118 3548 3152
rect 3582 3118 3620 3152
rect 3654 3118 3692 3152
rect 3726 3118 3794 3152
rect 2920 3112 3794 3118
tri 3834 3112 3878 3156 se
rect 3878 3112 3960 3156
tri 2920 3087 2945 3112 nw
tri 3809 3087 3834 3112 se
rect 3834 3087 3960 3112
tri 3806 3084 3809 3087 se
rect 3809 3084 3960 3087
rect 1753 3032 1931 3045
rect 1753 2980 1784 3032
rect 1836 2980 1848 3032
rect 1900 2980 1931 3032
rect 1753 2967 1931 2980
rect 1753 2915 1784 2967
rect 1836 2915 1848 2967
rect 1900 2915 1931 2967
rect 1753 2902 1931 2915
rect 1753 2850 1784 2902
rect 1836 2850 1848 2902
rect 1900 2850 1931 2902
tri 2948 3065 2967 3084 se
rect 2967 3065 3960 3084
rect 2948 3040 3960 3065
rect 2948 3010 3854 3040
rect 2948 2894 2954 3010
rect 3070 2968 3854 3010
tri 3854 2968 3926 3040 nw
rect 3070 2894 3076 2968
tri 3076 2943 3101 2968 nw
rect 1753 2837 1931 2850
rect 1753 2785 1784 2837
rect 1836 2785 1848 2837
rect 1900 2785 1931 2837
rect 1753 2772 1931 2785
rect 1753 2720 1784 2772
rect 1836 2720 1848 2772
rect 1900 2720 1931 2772
rect 1753 2714 1931 2720
rect 1518 2415 1544 2437
rect 998 2198 1130 2204
rect 998 2146 1006 2198
rect 1058 2146 1070 2198
rect 1122 2146 1130 2198
rect 998 2099 1130 2146
rect 1932 2198 2064 2204
rect 1932 2146 1940 2198
rect 1992 2146 2004 2198
rect 2056 2146 2064 2198
rect 998 2047 1006 2099
rect 1058 2047 1070 2099
rect 1122 2047 1130 2099
rect 998 2041 1130 2047
rect 1131 2132 1309 2138
rect 1131 2080 1162 2132
rect 1214 2080 1226 2132
rect 1278 2080 1309 2132
rect 1131 2067 1309 2080
tri 964 1976 1021 2033 sw
rect 1131 2015 1162 2067
rect 1214 2015 1226 2067
rect 1278 2015 1309 2067
rect 1131 2002 1309 2015
rect 948 1944 1021 1976
tri 1021 1944 1053 1976 sw
rect 1131 1950 1162 2002
rect 1214 1950 1226 2002
rect 1278 1950 1309 2002
rect 1131 1944 1309 1950
rect 1753 2132 1931 2138
rect 1753 2080 1784 2132
rect 1836 2080 1848 2132
rect 1900 2080 1931 2132
rect 1753 2067 1931 2080
rect 1753 2015 1784 2067
rect 1836 2015 1848 2067
rect 1900 2015 1931 2067
rect 1932 2099 2064 2146
rect 1932 2047 1940 2099
rect 1992 2047 2004 2099
rect 2056 2047 2064 2099
rect 1932 2041 2064 2047
rect 1753 2002 1931 2015
rect 1753 1950 1784 2002
rect 1836 1950 1848 2002
rect 1900 1950 1931 2002
rect 1753 1944 1931 1950
rect 2108 1944 2114 2892
rect 2230 1944 2236 2892
rect 2948 2861 3076 2894
tri 3076 2861 3110 2895 sw
rect 2948 2855 3768 2861
rect 2948 2675 2954 2855
rect 3070 2675 3084 2855
rect 3200 2675 3524 2855
rect 2948 2669 3768 2675
rect 2839 2404 2865 2453
rect 2281 2179 2483 2203
rect 2281 2127 2287 2179
rect 2339 2127 2356 2179
rect 2408 2127 2425 2179
rect 2477 2127 2483 2179
rect 2281 2115 2483 2127
rect 2281 2063 2287 2115
rect 2339 2063 2356 2115
rect 2408 2063 2425 2115
rect 2477 2063 2483 2115
rect 2281 2039 2483 2063
rect 2488 2132 2628 2138
rect 2488 2080 2500 2132
rect 2552 2080 2564 2132
rect 2616 2080 2628 2132
rect 2488 2067 2628 2080
rect 2488 2015 2500 2067
rect 2552 2015 2564 2067
rect 2616 2015 2628 2067
rect 2488 2002 2628 2015
rect 2488 1950 2500 2002
rect 2552 1950 2564 2002
rect 2616 1950 2628 2002
rect 2488 1944 2628 1950
rect 895 1929 1053 1944
tri 1053 1929 1068 1944 sw
tri 838 1872 895 1929 ne
rect 895 1902 1068 1929
tri 1068 1902 1095 1929 sw
rect 895 1847 1095 1902
rect 647 1503 827 1509
rect 647 1381 827 1387
rect 1977 1503 2157 1509
rect 1977 1381 2157 1387
rect 2948 1353 3076 2669
tri 3076 2642 3103 2669 nw
rect 3271 2476 3278 2592
rect 3394 2557 3524 2592
tri 3524 2557 3559 2592 sw
rect 3394 2476 3971 2557
rect 3271 2439 3971 2476
rect 3106 2405 3508 2411
rect 3106 2353 3122 2405
rect 3174 2353 3186 2405
rect 3238 2353 3250 2405
rect 3302 2353 3314 2405
rect 3366 2353 3508 2405
rect 3106 2291 3508 2353
rect 3106 2239 3122 2291
rect 3174 2239 3186 2291
rect 3238 2239 3250 2291
rect 3302 2239 3314 2291
rect 3366 2239 3508 2291
rect 3106 2233 3508 2239
rect 3524 1727 3962 1739
rect 3768 1547 3962 1727
rect 3524 1537 3962 1547
rect 439 1237 445 1353
rect 561 1237 567 1353
rect 1167 1237 1173 1353
rect 1289 1237 1295 1353
rect 1780 1237 1786 1353
rect 1902 1237 1908 1353
rect 2499 1237 2505 1353
rect 2621 1237 2627 1353
rect 2948 1237 2954 1353
rect 3070 1237 3076 1353
rect 3524 894 4014 923
rect 3768 778 4014 894
rect 3524 741 4014 778
rect 276 227 282 343
rect 590 227 596 343
rect 1468 227 1474 343
rect 1590 227 1596 343
rect 2230 227 2236 343
rect 2416 227 2422 343
rect 2467 227 2473 343
rect 2781 227 2787 343
rect 3106 -329 3508 -37
<< via1 >>
rect 282 4510 590 4626
rect 1474 4510 1590 4626
rect 2236 4606 2416 4626
rect 2236 4572 2238 4606
rect 2238 4572 2272 4606
rect 2272 4572 2310 4606
rect 2310 4572 2344 4606
rect 2344 4572 2382 4606
rect 2382 4572 2416 4606
rect 2236 4510 2416 4572
rect 2461 4510 2705 4626
rect 446 4066 562 4182
rect 1164 4066 1280 4182
rect 1786 4066 1902 4182
rect 2501 4066 2617 4182
rect 2959 4152 3075 4182
rect 2959 4118 3074 4152
rect 3074 4118 3075 4152
rect 2959 4080 3075 4118
rect 2959 4066 3074 4080
rect 3074 4066 3075 4080
rect 645 3916 825 4032
rect 1977 3916 2157 4032
rect 446 3766 562 3882
rect 1165 3766 1281 3882
rect 1781 3766 1897 3882
rect 2501 3766 2617 3882
rect 905 2924 1085 3616
rect 1162 3110 1278 3610
rect 1162 3045 1214 3097
rect 1226 3045 1278 3097
rect 1162 2980 1214 3032
rect 1226 2980 1278 3032
rect 832 1944 948 2892
rect 1162 2915 1214 2967
rect 1226 2915 1278 2967
rect 1162 2850 1214 2902
rect 1226 2850 1278 2902
rect 1162 2785 1214 2837
rect 1226 2785 1278 2837
rect 1162 2720 1214 2772
rect 1226 2720 1278 2772
rect 1784 3110 1900 3610
rect 2954 3247 3070 3875
rect 3181 4063 3233 4072
rect 3181 4029 3190 4063
rect 3190 4029 3224 4063
rect 3224 4029 3233 4063
rect 3181 4020 3233 4029
rect 3181 3991 3233 4008
rect 3181 3957 3190 3991
rect 3190 3957 3224 3991
rect 3224 3957 3233 3991
rect 3437 4076 3489 4080
rect 3437 4042 3446 4076
rect 3446 4042 3480 4076
rect 3480 4042 3489 4076
rect 3437 4028 3489 4042
rect 3437 4004 3489 4016
rect 3437 3970 3446 4004
rect 3446 3970 3480 4004
rect 3480 3970 3489 4004
rect 3437 3964 3489 3970
rect 3556 4064 3562 4080
rect 3562 4064 3596 4080
rect 3596 4064 3608 4080
rect 3556 4028 3608 4064
rect 3556 3992 3562 4016
rect 3562 3992 3596 4016
rect 3596 3992 3608 4016
rect 3556 3964 3608 3992
rect 3716 4139 3748 4153
rect 3748 4139 3768 4153
rect 3716 4101 3768 4139
rect 3716 4067 3748 4089
rect 3748 4067 3768 4089
rect 3716 4037 3768 4067
rect 3716 3995 3748 4025
rect 3748 3995 3768 4025
rect 3716 3973 3768 3995
rect 3181 3956 3233 3957
rect 3181 3919 3233 3944
rect 3181 3892 3190 3919
rect 3190 3892 3224 3919
rect 3224 3892 3233 3919
rect 3181 3847 3233 3880
rect 3181 3828 3190 3847
rect 3190 3828 3224 3847
rect 3224 3828 3233 3847
rect 3181 3813 3190 3816
rect 3190 3813 3224 3816
rect 3224 3813 3233 3816
rect 3181 3775 3233 3813
rect 3181 3764 3190 3775
rect 3190 3764 3224 3775
rect 3224 3764 3233 3775
rect 3181 3741 3190 3752
rect 3190 3741 3224 3752
rect 3224 3741 3233 3752
rect 3181 3703 3233 3741
rect 3181 3700 3190 3703
rect 3190 3700 3224 3703
rect 3224 3700 3233 3703
rect 3437 3797 3489 3811
rect 3437 3763 3446 3797
rect 3446 3763 3480 3797
rect 3480 3763 3489 3797
rect 3437 3759 3489 3763
rect 3437 3725 3489 3747
rect 3437 3695 3446 3725
rect 3446 3695 3480 3725
rect 3480 3695 3489 3725
rect 3437 3653 3489 3683
rect 3437 3631 3446 3653
rect 3446 3631 3480 3653
rect 3480 3631 3489 3653
rect 3556 3804 3562 3838
rect 3562 3804 3596 3838
rect 3596 3804 3608 3838
rect 3556 3786 3608 3804
rect 3556 3766 3608 3774
rect 3556 3732 3562 3766
rect 3562 3732 3596 3766
rect 3596 3732 3608 3766
rect 3556 3722 3608 3732
rect 3556 3694 3608 3710
rect 3556 3660 3562 3694
rect 3562 3660 3596 3694
rect 3596 3660 3608 3694
rect 3556 3658 3608 3660
rect 3716 3838 3768 3839
rect 3716 3804 3748 3838
rect 3748 3804 3768 3838
rect 3716 3787 3768 3804
rect 3716 3766 3768 3775
rect 3716 3732 3748 3766
rect 3748 3732 3768 3766
rect 3716 3723 3768 3732
rect 3716 3694 3768 3711
rect 3716 3660 3748 3694
rect 3748 3660 3768 3694
rect 3716 3659 3768 3660
rect 3437 3581 3489 3619
rect 3437 3567 3446 3581
rect 3446 3567 3480 3581
rect 3480 3567 3489 3581
rect 3437 3547 3446 3555
rect 3446 3547 3480 3555
rect 3480 3547 3489 3555
rect 3437 3503 3489 3547
rect 3556 3520 3608 3533
rect 3556 3486 3562 3520
rect 3562 3486 3596 3520
rect 3596 3486 3608 3520
rect 3556 3481 3608 3486
rect 3556 3448 3608 3469
rect 3278 3420 3330 3429
rect 3278 3386 3283 3420
rect 3283 3386 3317 3420
rect 3317 3386 3330 3420
rect 3278 3377 3330 3386
rect 3342 3420 3394 3429
rect 3342 3386 3355 3420
rect 3355 3386 3389 3420
rect 3389 3386 3394 3420
rect 3342 3377 3394 3386
rect 3556 3417 3562 3448
rect 3562 3417 3596 3448
rect 3596 3417 3608 3448
rect 3556 3376 3608 3405
rect 3556 3353 3562 3376
rect 3562 3353 3596 3376
rect 3596 3353 3608 3376
rect 3716 3508 3768 3527
rect 3716 3475 3748 3508
rect 3748 3475 3768 3508
rect 3716 3436 3768 3463
rect 3716 3411 3748 3436
rect 3748 3411 3768 3436
rect 3716 3364 3768 3399
rect 3716 3347 3748 3364
rect 3748 3347 3768 3364
rect 3716 3330 3748 3335
rect 3748 3330 3768 3335
rect 3716 3292 3768 3330
rect 3716 3283 3748 3292
rect 3748 3283 3768 3292
rect 3716 3258 3748 3271
rect 3748 3258 3768 3271
rect 3716 3220 3768 3258
rect 3716 3219 3748 3220
rect 3748 3219 3768 3220
rect 3716 3186 3748 3207
rect 3748 3186 3768 3207
rect 1784 3045 1836 3097
rect 1848 3045 1900 3097
rect 3716 3155 3768 3186
rect 1784 2980 1836 3032
rect 1848 2980 1900 3032
rect 1784 2915 1836 2967
rect 1848 2915 1900 2967
rect 1784 2850 1836 2902
rect 1848 2850 1900 2902
rect 2954 2894 3070 3010
rect 1784 2785 1836 2837
rect 1848 2785 1900 2837
rect 1784 2720 1836 2772
rect 1848 2720 1900 2772
rect 1006 2146 1058 2198
rect 1070 2146 1122 2198
rect 1940 2146 1992 2198
rect 2004 2146 2056 2198
rect 1006 2047 1058 2099
rect 1070 2047 1122 2099
rect 1162 2080 1214 2132
rect 1226 2080 1278 2132
rect 1162 2015 1214 2067
rect 1226 2015 1278 2067
rect 1162 1950 1214 2002
rect 1226 1950 1278 2002
rect 1784 2080 1836 2132
rect 1848 2080 1900 2132
rect 1784 2015 1836 2067
rect 1848 2015 1900 2067
rect 1940 2047 1992 2099
rect 2004 2047 2056 2099
rect 1784 1950 1836 2002
rect 1848 1950 1900 2002
rect 2114 1944 2230 2892
rect 2954 2675 3070 2855
rect 3084 2675 3200 2855
rect 3524 2675 3768 2855
rect 2287 2127 2339 2179
rect 2356 2127 2408 2179
rect 2425 2127 2477 2179
rect 2287 2063 2339 2115
rect 2356 2063 2408 2115
rect 2425 2063 2477 2115
rect 2500 2080 2552 2132
rect 2564 2080 2616 2132
rect 2500 2015 2552 2067
rect 2564 2015 2616 2067
rect 2500 1950 2552 2002
rect 2564 1950 2616 2002
rect 647 1387 827 1503
rect 1977 1387 2157 1503
rect 3278 2476 3394 2592
rect 3122 2353 3174 2405
rect 3186 2353 3238 2405
rect 3250 2353 3302 2405
rect 3314 2353 3366 2405
rect 3122 2239 3174 2291
rect 3186 2239 3238 2291
rect 3250 2239 3302 2291
rect 3314 2239 3366 2291
rect 3524 1547 3768 1727
rect 445 1237 561 1353
rect 1173 1237 1289 1353
rect 1786 1237 1902 1353
rect 2505 1237 2621 1353
rect 2954 1237 3070 1353
rect 3524 778 3768 894
rect 282 227 590 343
rect 1474 227 1590 343
rect 2236 280 2416 343
rect 2236 246 2238 280
rect 2238 246 2272 280
rect 2272 246 2310 280
rect 2310 246 2344 280
rect 2344 246 2382 280
rect 2382 246 2416 280
rect 2236 227 2416 246
rect 2473 227 2781 343
<< metal2 >>
rect 276 4510 282 4626
rect 590 4510 1474 4626
rect 1590 4510 2236 4626
rect 2416 4510 2461 4626
rect 2705 4510 2711 4626
rect 440 4066 446 4182
rect 562 4066 1164 4182
rect 1280 4066 1786 4182
rect 1902 4066 2501 4182
rect 2617 4066 2959 4182
rect 3075 4066 3081 4182
rect 3716 4153 3768 4159
rect 3716 4089 3768 4101
rect 3437 4080 3489 4086
tri 3177 4072 3181 4076 se
rect 3181 4072 3233 4078
tri 3171 4066 3177 4072 se
rect 3177 4066 3181 4072
tri 3143 4038 3171 4066 se
rect 3171 4038 3181 4066
rect 148 4032 3181 4038
rect 148 3916 645 4032
rect 825 3916 1977 4032
rect 2157 4020 3181 4032
rect 2157 4008 3233 4020
rect 2157 3956 3181 4008
rect 2157 3944 3233 3956
rect 2157 3916 3181 3944
rect 148 3910 3181 3916
rect 148 3892 410 3910
tri 410 3892 428 3910 nw
tri 3143 3892 3161 3910 ne
rect 3161 3892 3181 3910
rect 148 1944 403 3892
tri 403 3885 410 3892 nw
tri 3161 3885 3168 3892 ne
rect 3168 3885 3233 3892
tri 3168 3882 3171 3885 ne
rect 3171 3882 3233 3885
rect 440 3766 446 3882
rect 562 3766 1165 3882
rect 1281 3766 1781 3882
rect 1897 3766 2501 3882
rect 2617 3875 3076 3882
tri 3171 3880 3173 3882 ne
rect 3173 3880 3233 3882
rect 2617 3766 2954 3875
tri 2922 3740 2948 3766 ne
rect 826 2924 905 3616
rect 1085 3610 2667 3616
rect 1085 3110 1162 3610
rect 1278 3110 1784 3610
rect 1900 3110 2667 3610
rect 1085 3097 2667 3110
rect 1085 3045 1162 3097
rect 1214 3045 1226 3097
rect 1278 3045 1784 3097
rect 1836 3045 1848 3097
rect 1900 3045 2667 3097
rect 1085 3032 2667 3045
rect 1085 2980 1162 3032
rect 1214 2980 1226 3032
rect 1278 2980 1784 3032
rect 1836 2980 1848 3032
rect 1900 2980 2667 3032
rect 1085 2967 2667 2980
rect 1085 2924 1162 2967
rect 826 2915 1162 2924
rect 1214 2915 1226 2967
rect 1278 2915 1784 2967
rect 1836 2915 1848 2967
rect 1900 2915 2667 2967
rect 826 2902 2667 2915
rect 826 2892 1162 2902
tri 403 1944 496 2037 sw
rect 826 1944 832 2892
rect 948 2850 1162 2892
rect 1214 2850 1226 2902
rect 1278 2850 1784 2902
rect 1836 2850 1848 2902
rect 1900 2892 2667 2902
rect 1900 2850 2114 2892
rect 948 2837 2114 2850
rect 948 2785 1162 2837
rect 1214 2785 1226 2837
rect 1278 2785 1784 2837
rect 1836 2785 1848 2837
rect 1900 2785 2114 2837
rect 948 2772 2114 2785
rect 948 2720 1162 2772
rect 1214 2720 1226 2772
rect 1278 2720 1784 2772
rect 1836 2720 1848 2772
rect 1900 2720 2114 2772
rect 948 2198 2114 2720
rect 948 2146 1006 2198
rect 1058 2146 1070 2198
rect 1122 2146 1940 2198
rect 1992 2146 2004 2198
rect 2056 2146 2114 2198
rect 948 2132 2114 2146
rect 948 2099 1162 2132
rect 948 2047 1006 2099
rect 1058 2047 1070 2099
rect 1122 2080 1162 2099
rect 1214 2080 1226 2132
rect 1278 2080 1784 2132
rect 1836 2080 1848 2132
rect 1900 2099 2114 2132
rect 1900 2080 1940 2099
rect 1122 2067 1940 2080
rect 1122 2047 1162 2067
rect 948 2015 1162 2047
rect 1214 2015 1226 2067
rect 1278 2015 1784 2067
rect 1836 2015 1848 2067
rect 1900 2047 1940 2067
rect 1992 2047 2004 2099
rect 2056 2047 2114 2099
rect 1900 2015 2114 2047
rect 948 2002 2114 2015
rect 948 1950 1162 2002
rect 1214 1950 1226 2002
rect 1278 1950 1784 2002
rect 1836 1950 1848 2002
rect 1900 1950 2114 2002
rect 948 1944 2114 1950
rect 2230 2252 2667 2892
rect 2948 3247 2954 3766
rect 3070 3247 3076 3875
tri 3173 3872 3181 3880 ne
rect 3181 3816 3233 3828
rect 3181 3752 3233 3764
rect 3181 3694 3233 3700
rect 3437 4016 3489 4028
rect 3437 3811 3489 3964
rect 3437 3747 3489 3759
rect 3437 3683 3489 3695
rect 3437 3619 3489 3631
rect 3437 3555 3489 3567
rect 2948 3010 3076 3247
rect 2948 2894 2954 3010
rect 3070 2894 3076 3010
rect 2948 2861 3076 2894
rect 3272 3377 3278 3429
rect 3330 3377 3342 3429
rect 3394 3377 3400 3429
rect 2948 2855 3200 2861
rect 2948 2675 2954 2855
rect 3070 2675 3084 2855
rect 2948 2669 3200 2675
rect 2948 2252 3066 2669
rect 3272 2592 3400 3377
rect 3437 2769 3489 3503
rect 3556 4080 3608 4086
rect 3556 4016 3608 4028
rect 3556 3838 3608 3964
rect 3556 3774 3608 3786
rect 3556 3710 3608 3722
rect 3556 3533 3608 3658
rect 3556 3469 3608 3481
rect 3556 3405 3608 3417
rect 3556 3347 3608 3353
rect 3716 4025 3768 4037
rect 3716 3839 3768 3973
rect 3716 3775 3768 3787
rect 3716 3711 3768 3723
rect 3716 3527 3768 3659
rect 3716 3463 3768 3475
rect 3716 3399 3768 3411
rect 3716 3335 3768 3347
rect 3716 3271 3768 3283
rect 3716 3207 3768 3219
rect 3716 3149 3768 3155
rect 3524 2855 3768 2861
tri 3489 2769 3496 2776 sw
rect 3437 2754 3496 2769
tri 3437 2747 3444 2754 ne
rect 3272 2476 3278 2592
rect 3394 2476 3400 2592
rect 2230 2179 3066 2252
rect 2230 2127 2287 2179
rect 2339 2127 2356 2179
rect 2408 2127 2425 2179
rect 2477 2132 3066 2179
rect 2477 2127 2500 2132
rect 2230 2115 2500 2127
rect 2230 2063 2287 2115
rect 2339 2063 2356 2115
rect 2408 2063 2425 2115
rect 2477 2080 2500 2115
rect 2552 2080 2564 2132
rect 2616 2080 3066 2132
rect 2477 2067 3066 2080
rect 2477 2063 2500 2067
rect 2230 2015 2500 2063
rect 2552 2015 2564 2067
rect 2616 2060 3066 2067
rect 3106 2405 3412 2411
rect 3106 2353 3122 2405
rect 3174 2353 3186 2405
rect 3238 2353 3250 2405
rect 3302 2353 3314 2405
rect 3366 2353 3412 2405
rect 3106 2291 3412 2353
rect 3106 2239 3122 2291
rect 3174 2239 3186 2291
rect 3238 2239 3250 2291
rect 3302 2239 3314 2291
rect 3366 2239 3412 2291
rect 2616 2034 3025 2060
tri 3025 2034 3051 2060 nw
rect 2616 2015 2960 2034
rect 2230 2002 2960 2015
rect 2230 1950 2500 2002
rect 2552 1950 2564 2002
rect 2616 1969 2960 2002
tri 2960 1969 3025 2034 nw
tri 3041 1969 3106 2034 se
rect 3106 1969 3412 2239
rect 2616 1950 2935 1969
rect 2230 1944 2935 1950
tri 2935 1944 2960 1969 nw
tri 3016 1944 3041 1969 se
rect 3041 1944 3412 1969
rect 148 1888 496 1944
tri 496 1888 552 1944 sw
tri 2960 1888 3016 1944 se
rect 3016 1888 3412 1944
rect 148 1571 3412 1888
rect 148 1547 3388 1571
tri 3388 1547 3412 1571 nw
rect 148 1537 3378 1547
tri 3378 1537 3388 1547 nw
tri 3434 1537 3444 1547 se
rect 3444 1537 3496 2754
tri 3406 1509 3434 1537 se
rect 3434 1509 3496 1537
rect 647 1503 3496 1509
rect 827 1387 1977 1503
rect 2157 1387 3496 1503
rect 647 1381 3496 1387
rect 3524 1727 3768 2675
rect 437 1237 445 1353
rect 561 1237 1173 1353
rect 1289 1237 1786 1353
rect 1902 1237 2505 1353
rect 2621 1237 2954 1353
rect 3070 1237 3076 1353
rect 3524 894 3768 1547
rect 3524 772 3768 778
rect 276 227 282 343
rect 590 227 1474 343
rect 1590 227 2236 343
rect 2416 227 2473 343
rect 2781 227 2787 343
use sky130_fd_io__res250only_small  sky130_fd_io__res250only_small_0
timestamp 1681267127
transform 0 -1 3509 1 0 -37
box 0 0 2270 404
use sky130_fd_io__signal_5_sym_hv_local_5term  sky130_fd_io__signal_5_sym_hv_local_5term_0
timestamp 1681267127
transform 1 0 1395 0 1 138
box 0 0 1591 2424
use sky130_fd_io__signal_5_sym_hv_local_5term  sky130_fd_io__signal_5_sym_hv_local_5term_1
timestamp 1681267127
transform -1 0 1667 0 1 138
box 0 0 1591 2424
use sky130_fd_io__signal_5_sym_hv_local_5term  sky130_fd_io__signal_5_sym_hv_local_5term_2
timestamp 1681267127
transform 1 0 1395 0 -1 4714
box 0 0 1591 2424
use sky130_fd_io__signal_5_sym_hv_local_5term  sky130_fd_io__signal_5_sym_hv_local_5term_3
timestamp 1681267127
transform -1 0 1667 0 -1 4714
box 0 0 1591 2424
use sky130_fd_pr__nfet_01v8__example_55959141808555  sky130_fd_pr__nfet_01v8__example_55959141808555_0
timestamp 1681267127
transform -1 0 3435 0 -1 4062
box -1 0 201 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_0
timestamp 1681267127
transform 0 1 3446 -1 0 4076
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_1
timestamp 1681267127
transform 1 0 3283 0 -1 3420
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_0
timestamp 1681267127
transform 0 -1 3782 -1 0 3838
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_1
timestamp 1681267127
transform 0 -1 3596 1 0 3660
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_2
timestamp 1681267127
transform 0 -1 3596 1 0 3342
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_3
timestamp 1681267127
transform 0 -1 3596 -1 0 4170
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808127  sky130_fd_pr__via_l1m1__example_55959141808127_0
timestamp 1681267127
transform 0 1 3446 1 0 3547
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808127  sky130_fd_pr__via_l1m1__example_55959141808127_1
timestamp 1681267127
transform 0 -1 3782 1 0 3995
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808128  sky130_fd_pr__via_l1m1__example_55959141808128_0
timestamp 1681267127
transform 0 1 2238 -1 0 280
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808128  sky130_fd_pr__via_l1m1__example_55959141808128_1
timestamp 1681267127
transform 0 1 2238 -1 0 4606
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808290  sky130_fd_pr__via_l1m1__example_55959141808290_0
timestamp 1681267127
transform 0 1 3190 1 0 3525
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808326  sky130_fd_pr__via_l1m1__example_55959141808326_0
timestamp 1681267127
transform -1 0 3726 0 -1 3152
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808326  sky130_fd_pr__via_l1m1__example_55959141808326_1
timestamp 1681267127
transform 1 0 2975 0 -1 4356
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808372  sky130_fd_pr__via_l1m1__example_55959141808372_0
timestamp 1681267127
transform 1 0 3169 0 -1 4170
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808372  sky130_fd_pr__via_l1m1__example_55959141808372_1
timestamp 1681267127
transform 0 -1 3782 1 0 3186
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808400  sky130_fd_pr__via_l1m1__example_55959141808400_0
timestamp 1681267127
transform 0 -1 3108 1 0 3326
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808259  sky130_fd_pr__via_m1m2__example_55959141808259_0
timestamp 1681267127
transform 0 1 3437 1 0 3497
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_0
timestamp 1681267127
transform 0 1 3437 -1 0 4086
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_1
timestamp 1681267127
transform 0 1 3556 -1 0 4086
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_2
timestamp 1681267127
transform -1 0 3400 0 -1 3429
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808261  sky130_fd_pr__via_m1m2__example_55959141808261_0
timestamp 1681267127
transform 0 -1 3768 1 0 3967
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808261  sky130_fd_pr__via_m1m2__example_55959141808261_1
timestamp 1681267127
transform 0 -1 3768 1 0 3653
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808261  sky130_fd_pr__via_m1m2__example_55959141808261_2
timestamp 1681267127
transform 0 1 3556 -1 0 3539
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808261  sky130_fd_pr__via_m1m2__example_55959141808261_3
timestamp 1681267127
transform 0 1 3556 -1 0 3844
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808350  sky130_fd_pr__via_m1m2__example_55959141808350_0
timestamp 1681267127
transform 1 0 2948 0 -1 3010
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808350  sky130_fd_pr__via_m1m2__example_55959141808350_1
timestamp 1681267127
transform -1 0 3400 0 -1 2592
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808350  sky130_fd_pr__via_m1m2__example_55959141808350_2
timestamp 1681267127
transform 1 0 1468 0 1 227
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808350  sky130_fd_pr__via_m1m2__example_55959141808350_3
timestamp 1681267127
transform 1 0 1468 0 1 4510
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808350  sky130_fd_pr__via_m1m2__example_55959141808350_4
timestamp 1681267127
transform -1 0 2627 0 -1 1353
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808350  sky130_fd_pr__via_m1m2__example_55959141808350_5
timestamp 1681267127
transform 1 0 439 0 -1 1353
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808350  sky130_fd_pr__via_m1m2__example_55959141808350_6
timestamp 1681267127
transform 1 0 440 0 -1 4182
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808350  sky130_fd_pr__via_m1m2__example_55959141808350_7
timestamp 1681267127
transform 1 0 1158 0 -1 4182
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808350  sky130_fd_pr__via_m1m2__example_55959141808350_8
timestamp 1681267127
transform 1 0 1780 0 -1 4182
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808350  sky130_fd_pr__via_m1m2__example_55959141808350_9
timestamp 1681267127
transform 1 0 2495 0 -1 3882
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808350  sky130_fd_pr__via_m1m2__example_55959141808350_10
timestamp 1681267127
transform 1 0 440 0 -1 3882
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808350  sky130_fd_pr__via_m1m2__example_55959141808350_11
timestamp 1681267127
transform 1 0 2495 0 1 4066
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808350  sky130_fd_pr__via_m1m2__example_55959141808350_12
timestamp 1681267127
transform 1 0 2953 0 1 4066
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808350  sky130_fd_pr__via_m1m2__example_55959141808350_13
timestamp 1681267127
transform 1 0 1780 0 -1 1353
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808350  sky130_fd_pr__via_m1m2__example_55959141808350_14
timestamp 1681267127
transform -1 0 1295 0 -1 1353
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808350  sky130_fd_pr__via_m1m2__example_55959141808350_15
timestamp 1681267127
transform 1 0 1159 0 -1 3882
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808350  sky130_fd_pr__via_m1m2__example_55959141808350_16
timestamp 1681267127
transform 1 0 2948 0 -1 1353
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808350  sky130_fd_pr__via_m1m2__example_55959141808350_17
timestamp 1681267127
transform 1 0 1775 0 -1 3882
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808402  sky130_fd_pr__via_m1m2__example_55959141808402_0
timestamp 1681267127
transform 0 1 647 1 0 1381
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808402  sky130_fd_pr__via_m1m2__example_55959141808402_1
timestamp 1681267127
transform 0 1 645 1 0 3910
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808402  sky130_fd_pr__via_m1m2__example_55959141808402_2
timestamp 1681267127
transform 0 1 1977 1 0 1381
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808402  sky130_fd_pr__via_m1m2__example_55959141808402_3
timestamp 1681267127
transform 0 1 1977 1 0 3910
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808551  sky130_fd_pr__via_m1m2__example_55959141808551_0
timestamp 1681267127
transform -1 0 2711 0 1 4510
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808552  sky130_fd_pr__via_m1m2__example_55959141808552_0
timestamp 1681267127
transform 1 0 2230 0 1 4510
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808552  sky130_fd_pr__via_m1m2__example_55959141808552_1
timestamp 1681267127
transform 0 1 3084 -1 0 2861
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808552  sky130_fd_pr__via_m1m2__example_55959141808552_2
timestamp 1681267127
transform 1 0 2230 0 1 227
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808553  sky130_fd_pr__via_m1m2__example_55959141808553_0
timestamp 1681267127
transform 0 -1 3768 -1 0 3533
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808553  sky130_fd_pr__via_m1m2__example_55959141808553_1
timestamp 1681267127
transform 0 1 3181 -1 0 4078
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808554  sky130_fd_pr__via_m1m2__example_55959141808554_0
timestamp 1681267127
transform 1 0 2108 0 1 1944
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808554  sky130_fd_pr__via_m1m2__example_55959141808554_1
timestamp 1681267127
transform 1 0 826 0 1 1944
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808724  sky130_fd_pr__via_m1m2__example_55959141808724_0
timestamp 1681267127
transform -1 0 2787 0 1 227
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808724  sky130_fd_pr__via_m1m2__example_55959141808724_1
timestamp 1681267127
transform -1 0 596 0 1 227
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808724  sky130_fd_pr__via_m1m2__example_55959141808724_2
timestamp 1681267127
transform -1 0 596 0 1 4510
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808725  sky130_fd_pr__via_m1m2__example_55959141808725_0
timestamp 1681267127
transform 1 0 2948 0 1 3247
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808726  sky130_fd_pr__via_m1m2__example_55959141808726_0
timestamp 1681267127
transform 1 0 899 0 -1 3616
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808727  sky130_fd_pr__via_m1m2__example_55959141808727_0
timestamp 1681267127
transform 0 1 3524 -1 0 2861
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808727  sky130_fd_pr__via_m1m2__example_55959141808727_1
timestamp 1681267127
transform 0 1 3524 -1 0 1733
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808728  sky130_fd_pr__via_m1m2__example_55959141808728_0
timestamp 1681267127
transform 0 1 3524 -1 0 900
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808274  sky130_fd_pr__via_pol1__example_55959141808274_0
timestamp 1681267127
transform 0 1 3235 -1 0 3436
box 0 0 1 1
<< labels >>
flabel comment s 59 4554 59 4554 0 FreeSans 200 0 0 0 PAD
flabel metal2 s 1424 4525 1635 4597 0 FreeSans 200 0 0 0 VCC_IO
port 1 nsew
flabel metal1 s 3813 2472 3934 2523 0 FreeSans 200 0 0 0 VTRIP_SEL_H
port 3 nsew
flabel metal1 s 3952 1537 3962 1739 7 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel metal1 s 3975 3881 4014 3927 7 FreeSans 200 0 0 0 OUT_H
port 5 nsew
flabel metal1 s 3975 3571 4014 3617 7 FreeSans 200 0 0 0 OUT_VT
port 6 nsew
<< properties >>
string GDS_END 31287198
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 31261530
<< end >>
