magic
tech sky130A
magscale 1 2
timestamp 1681267127
<< nwell >>
rect -38 261 1510 582
<< pwell >>
rect 1 21 1471 203
rect 30 -17 64 21
<< locali >>
rect 27 149 70 325
rect 212 257 251 325
rect 543 309 777 343
rect 212 215 301 257
rect 582 177 621 309
rect 903 215 989 257
rect 1051 215 1208 257
rect 459 143 661 177
rect 459 93 493 143
rect 439 59 509 93
rect 627 93 661 143
rect 611 59 677 93
rect 1389 215 1455 323
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 35 459 405 493
rect 35 359 69 459
rect 103 391 169 425
rect 119 177 153 391
rect 203 359 237 459
rect 287 325 321 425
rect 371 359 405 459
rect 459 451 525 527
rect 627 451 693 527
rect 795 451 861 527
rect 895 417 929 493
rect 963 451 1035 527
rect 1075 417 1109 493
rect 1143 451 1209 527
rect 1319 417 1353 493
rect 439 383 1353 417
rect 439 325 477 383
rect 895 359 929 383
rect 1075 359 1109 383
rect 1319 359 1353 383
rect 1387 359 1454 527
rect 287 291 477 325
rect 371 215 541 249
rect 371 177 405 215
rect 830 291 1337 325
rect 830 249 864 291
rect 655 215 864 249
rect 119 143 405 177
rect 19 17 69 113
rect 119 93 153 143
rect 103 59 169 93
rect 203 17 237 109
rect 287 93 321 143
rect 271 59 337 93
rect 371 17 405 109
rect 543 17 577 109
rect 871 143 1201 177
rect 711 17 813 109
rect 871 93 905 143
rect 1135 129 1201 143
rect 855 59 921 93
rect 955 17 989 109
rect 1235 93 1269 177
rect 1303 165 1337 291
rect 1303 129 1369 165
rect 1403 100 1454 181
rect 1051 85 1269 93
rect 1387 85 1454 100
rect 1051 51 1454 85
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
<< metal1 >>
rect 0 561 1472 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 0 496 1472 527
rect 0 17 1472 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
rect 0 -48 1472 -17
<< labels >>
rlabel locali s 1389 215 1455 323 6 A1
port 1 nsew signal input
rlabel locali s 1051 215 1208 257 6 A2
port 2 nsew signal input
rlabel locali s 903 215 989 257 6 A3
port 3 nsew signal input
rlabel locali s 212 215 301 257 6 B1
port 4 nsew signal input
rlabel locali s 212 257 251 325 6 B1
port 4 nsew signal input
rlabel locali s 27 149 70 325 6 C1
port 5 nsew signal input
rlabel metal1 s 0 -48 1472 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 1 21 1471 203 6 VNB
port 7 nsew ground bidirectional
rlabel nwell s -38 261 1510 582 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 496 1472 592 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 611 59 677 93 6 X
port 10 nsew signal output
rlabel locali s 439 59 509 93 6 X
port 10 nsew signal output
rlabel locali s 627 93 661 143 6 X
port 10 nsew signal output
rlabel locali s 459 93 493 143 6 X
port 10 nsew signal output
rlabel locali s 459 143 661 177 6 X
port 10 nsew signal output
rlabel locali s 582 177 621 309 6 X
port 10 nsew signal output
rlabel locali s 543 309 777 343 6 X
port 10 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1472 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 3720592
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3708870
<< end >>
