magic
tech sky130A
magscale 1 2
timestamp 1681267127
<< nwell >>
rect -38 261 1050 582
<< pwell >>
rect 1 21 975 203
rect 30 -17 64 21
<< scnmos >>
rect 83 47 113 177
rect 167 47 197 177
rect 251 47 281 177
rect 335 47 365 177
rect 419 47 449 177
rect 503 47 533 177
rect 587 47 617 177
rect 671 47 701 177
rect 865 47 895 177
<< scpmoshvt >>
rect 83 297 113 497
rect 167 297 197 497
rect 251 297 281 497
rect 335 297 365 497
rect 419 297 449 497
rect 503 297 533 497
rect 587 297 617 497
rect 671 297 701 497
rect 865 297 895 497
<< ndiff >>
rect 27 163 83 177
rect 27 129 39 163
rect 73 129 83 163
rect 27 95 83 129
rect 27 61 39 95
rect 73 61 83 95
rect 27 47 83 61
rect 113 163 167 177
rect 113 129 123 163
rect 157 129 167 163
rect 113 95 167 129
rect 113 61 123 95
rect 157 61 167 95
rect 113 47 167 61
rect 197 95 251 177
rect 197 61 207 95
rect 241 61 251 95
rect 197 47 251 61
rect 281 163 335 177
rect 281 129 291 163
rect 325 129 335 163
rect 281 95 335 129
rect 281 61 291 95
rect 325 61 335 95
rect 281 47 335 61
rect 365 95 419 177
rect 365 61 375 95
rect 409 61 419 95
rect 365 47 419 61
rect 449 163 503 177
rect 449 129 459 163
rect 493 129 503 163
rect 449 95 503 129
rect 449 61 459 95
rect 493 61 503 95
rect 449 47 503 61
rect 533 95 587 177
rect 533 61 543 95
rect 577 61 587 95
rect 533 47 587 61
rect 617 163 671 177
rect 617 129 627 163
rect 661 129 671 163
rect 617 95 671 129
rect 617 61 627 95
rect 661 61 671 95
rect 617 47 671 61
rect 701 163 753 177
rect 701 129 711 163
rect 745 129 753 163
rect 701 95 753 129
rect 701 61 711 95
rect 745 61 753 95
rect 701 47 753 61
rect 809 163 865 177
rect 809 129 821 163
rect 855 129 865 163
rect 809 95 865 129
rect 809 61 821 95
rect 855 61 865 95
rect 809 47 865 61
rect 895 163 949 177
rect 895 129 905 163
rect 939 129 949 163
rect 895 95 949 129
rect 895 61 905 95
rect 939 61 949 95
rect 895 47 949 61
<< pdiff >>
rect 27 477 83 497
rect 27 443 39 477
rect 73 443 83 477
rect 27 409 83 443
rect 27 375 39 409
rect 73 375 83 409
rect 27 341 83 375
rect 27 307 39 341
rect 73 307 83 341
rect 27 297 83 307
rect 113 485 167 497
rect 113 451 123 485
rect 157 451 167 485
rect 113 417 167 451
rect 113 383 123 417
rect 157 383 167 417
rect 113 297 167 383
rect 197 477 251 497
rect 197 443 207 477
rect 241 443 251 477
rect 197 409 251 443
rect 197 375 207 409
rect 241 375 251 409
rect 197 341 251 375
rect 197 307 207 341
rect 241 307 251 341
rect 197 297 251 307
rect 281 485 335 497
rect 281 451 291 485
rect 325 451 335 485
rect 281 417 335 451
rect 281 383 291 417
rect 325 383 335 417
rect 281 297 335 383
rect 365 485 419 497
rect 365 451 375 485
rect 409 451 419 485
rect 365 417 419 451
rect 365 383 375 417
rect 409 383 419 417
rect 365 341 419 383
rect 365 307 375 341
rect 409 307 419 341
rect 365 297 419 307
rect 449 409 503 497
rect 449 375 459 409
rect 493 375 503 409
rect 449 341 503 375
rect 449 307 459 341
rect 493 307 503 341
rect 449 297 503 307
rect 533 489 587 497
rect 533 455 543 489
rect 577 455 587 489
rect 533 421 587 455
rect 533 387 543 421
rect 577 387 587 421
rect 533 297 587 387
rect 617 409 671 497
rect 617 375 627 409
rect 661 375 671 409
rect 617 341 671 375
rect 617 307 627 341
rect 661 307 671 341
rect 617 297 671 307
rect 701 485 757 497
rect 701 451 711 485
rect 745 451 757 485
rect 701 417 757 451
rect 701 383 711 417
rect 745 383 757 417
rect 701 349 757 383
rect 701 315 711 349
rect 745 315 757 349
rect 701 297 757 315
rect 811 485 865 497
rect 811 451 821 485
rect 855 451 865 485
rect 811 417 865 451
rect 811 383 821 417
rect 855 383 865 417
rect 811 349 865 383
rect 811 315 821 349
rect 855 315 865 349
rect 811 297 865 315
rect 895 485 951 497
rect 895 451 905 485
rect 939 451 951 485
rect 895 417 951 451
rect 895 383 905 417
rect 939 383 951 417
rect 895 349 951 383
rect 895 315 905 349
rect 939 315 951 349
rect 895 297 951 315
<< ndiffc >>
rect 39 129 73 163
rect 39 61 73 95
rect 123 129 157 163
rect 123 61 157 95
rect 207 61 241 95
rect 291 129 325 163
rect 291 61 325 95
rect 375 61 409 95
rect 459 129 493 163
rect 459 61 493 95
rect 543 61 577 95
rect 627 129 661 163
rect 627 61 661 95
rect 711 129 745 163
rect 711 61 745 95
rect 821 129 855 163
rect 821 61 855 95
rect 905 129 939 163
rect 905 61 939 95
<< pdiffc >>
rect 39 443 73 477
rect 39 375 73 409
rect 39 307 73 341
rect 123 451 157 485
rect 123 383 157 417
rect 207 443 241 477
rect 207 375 241 409
rect 207 307 241 341
rect 291 451 325 485
rect 291 383 325 417
rect 375 451 409 485
rect 375 383 409 417
rect 375 307 409 341
rect 459 375 493 409
rect 459 307 493 341
rect 543 455 577 489
rect 543 387 577 421
rect 627 375 661 409
rect 627 307 661 341
rect 711 451 745 485
rect 711 383 745 417
rect 711 315 745 349
rect 821 451 855 485
rect 821 383 855 417
rect 821 315 855 349
rect 905 451 939 485
rect 905 383 939 417
rect 905 315 939 349
<< poly >>
rect 83 249 365 265
rect 83 215 103 249
rect 137 215 171 249
rect 205 215 239 249
rect 273 215 307 249
rect 341 215 365 249
rect 83 199 365 215
rect 419 249 823 265
rect 419 215 575 249
rect 609 215 643 249
rect 677 215 711 249
rect 745 215 779 249
rect 813 215 823 249
rect 419 199 823 215
rect 865 249 955 265
rect 865 215 905 249
rect 939 215 955 249
rect 865 199 955 215
<< polycont >>
rect 103 215 137 249
rect 171 215 205 249
rect 239 215 273 249
rect 307 215 341 249
rect 575 215 609 249
rect 643 215 677 249
rect 711 215 745 249
rect 779 215 813 249
rect 905 215 939 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 17 477 73 493
rect 17 443 39 477
rect 17 409 73 443
rect 17 375 39 409
rect 17 341 73 375
rect 107 485 173 527
rect 107 451 123 485
rect 157 451 173 485
rect 107 417 173 451
rect 107 383 123 417
rect 157 383 173 417
rect 107 367 173 383
rect 207 477 241 493
rect 207 409 241 443
rect 17 307 39 341
rect 207 341 241 375
rect 275 485 325 527
rect 275 451 291 485
rect 275 417 325 451
rect 275 383 291 417
rect 275 367 325 383
rect 359 489 771 493
rect 359 485 543 489
rect 359 451 375 485
rect 409 459 543 485
rect 409 451 425 459
rect 359 417 425 451
rect 527 455 543 459
rect 577 485 771 489
rect 577 459 711 485
rect 577 455 593 459
rect 359 383 375 417
rect 409 383 425 417
rect 73 307 207 333
rect 359 341 425 383
rect 359 333 375 341
rect 241 307 375 333
rect 409 307 425 341
rect 17 291 425 307
rect 459 409 493 425
rect 527 421 593 455
rect 695 451 711 459
rect 745 451 771 485
rect 527 387 543 421
rect 577 387 593 421
rect 627 409 661 425
rect 459 349 493 375
rect 627 349 661 375
rect 459 341 661 349
rect 493 307 627 341
rect 695 417 771 451
rect 695 383 711 417
rect 745 383 771 417
rect 695 349 771 383
rect 695 315 711 349
rect 745 315 771 349
rect 805 485 871 493
rect 805 451 821 485
rect 855 451 871 485
rect 805 417 871 451
rect 805 383 821 417
rect 855 383 871 417
rect 805 349 871 383
rect 805 315 821 349
rect 855 315 871 349
rect 905 485 986 527
rect 939 451 986 485
rect 905 417 986 451
rect 939 383 986 417
rect 905 349 986 383
rect 939 315 986 349
rect 459 289 661 307
rect 72 249 360 255
rect 72 215 103 249
rect 137 215 171 249
rect 205 215 239 249
rect 273 215 307 249
rect 341 215 360 249
rect 459 181 525 289
rect 805 255 855 315
rect 905 299 986 315
rect 559 249 855 255
rect 559 215 575 249
rect 609 215 643 249
rect 677 215 711 249
rect 745 215 779 249
rect 813 215 855 249
rect 889 249 995 264
rect 889 215 905 249
rect 939 215 995 249
rect 17 163 73 181
rect 17 129 39 163
rect 17 95 73 129
rect 17 61 39 95
rect 17 17 73 61
rect 107 163 677 181
rect 107 129 123 163
rect 157 145 291 163
rect 157 129 173 145
rect 107 95 173 129
rect 275 129 291 145
rect 325 145 459 163
rect 325 129 341 145
rect 107 61 123 95
rect 157 61 173 95
rect 107 51 173 61
rect 207 95 241 111
rect 207 17 241 61
rect 275 95 341 129
rect 443 129 459 145
rect 493 145 627 163
rect 493 129 509 145
rect 275 61 291 95
rect 325 61 341 95
rect 275 51 341 61
rect 375 95 409 111
rect 375 17 409 61
rect 443 95 509 129
rect 611 129 627 145
rect 661 129 677 163
rect 443 61 459 95
rect 493 61 509 95
rect 443 51 509 61
rect 543 95 577 111
rect 543 17 577 61
rect 611 95 677 129
rect 611 61 627 95
rect 661 61 677 95
rect 611 51 677 61
rect 711 163 769 181
rect 745 129 769 163
rect 711 95 769 129
rect 745 61 769 95
rect 711 17 769 61
rect 805 163 855 215
rect 905 163 963 181
rect 805 129 821 163
rect 855 129 871 163
rect 805 95 871 129
rect 805 61 821 95
rect 855 61 871 95
rect 805 51 871 61
rect 939 129 963 163
rect 905 95 963 129
rect 939 61 963 95
rect 905 17 963 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
<< metal1 >>
rect 0 561 1012 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 0 496 1012 527
rect 0 17 1012 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
rect 0 -48 1012 -17
<< labels >>
flabel locali s 950 221 984 255 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 582 289 616 323 0 FreeSans 400 0 0 0 X
port 7 nsew signal output
flabel locali s 122 221 156 255 0 FreeSans 200 0 0 0 SLEEP
port 2 nsew signal input
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 lpflow_isobufsrc_4
rlabel metal1 s 0 -48 1012 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1012 592 1 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1012 544
string GDS_END 2385496
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2376978
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 25.300 0.000 
<< end >>
