magic
tech sky130A
magscale 1 2
timestamp 1681267127
<< nwell >>
rect -38 261 2062 582
<< pwell >>
rect 1 21 2023 203
rect 29 -17 63 21
<< locali >>
rect 20 199 66 323
rect 118 199 195 323
rect 508 333 558 493
rect 676 333 742 493
rect 844 333 910 493
rect 1012 333 1078 493
rect 1348 333 1414 493
rect 1516 333 1582 493
rect 1684 333 1750 493
rect 1852 333 1918 493
rect 508 289 1918 333
rect 740 181 798 289
rect 1224 215 1582 255
rect 1684 215 2003 255
rect 508 131 798 181
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 17 396 74 488
rect 108 439 153 527
rect 187 430 359 493
rect 17 357 291 396
rect 229 161 291 357
rect 17 127 291 161
rect 325 261 359 430
rect 440 299 474 527
rect 592 367 642 527
rect 776 367 810 527
rect 944 367 978 527
rect 1122 367 1308 527
rect 1448 367 1482 527
rect 1616 367 1650 527
rect 1784 367 1818 527
rect 1952 289 2007 527
rect 325 215 442 261
rect 508 215 657 249
rect 17 51 69 127
rect 325 93 359 215
rect 832 215 1078 255
rect 103 17 169 93
rect 203 51 359 93
rect 440 97 474 181
rect 844 147 1230 181
rect 844 131 1078 147
rect 1196 97 1230 147
rect 1264 131 2007 181
rect 440 51 1162 97
rect 1196 51 1582 97
rect 1684 17 1750 97
rect 1852 17 1918 97
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
<< metal1 >>
rect 0 561 2024 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 0 496 2024 527
rect 0 17 2024 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
rect 0 -48 2024 -17
<< obsm1 >>
rect 384 252 442 261
rect 844 252 902 261
rect 384 224 902 252
rect 384 215 442 224
rect 844 215 902 224
<< labels >>
rlabel locali s 20 199 66 323 6 A_N
port 1 nsew signal input
rlabel locali s 118 199 195 323 6 B_N
port 2 nsew signal input
rlabel locali s 1224 215 1582 255 6 C
port 3 nsew signal input
rlabel locali s 1684 215 2003 255 6 D
port 4 nsew signal input
rlabel metal1 s 0 -48 2024 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1 21 2023 203 6 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 2062 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 2024 592 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 508 131 798 181 6 Y
port 9 nsew signal output
rlabel locali s 740 181 798 289 6 Y
port 9 nsew signal output
rlabel locali s 508 289 1918 333 6 Y
port 9 nsew signal output
rlabel locali s 1852 333 1918 493 6 Y
port 9 nsew signal output
rlabel locali s 1684 333 1750 493 6 Y
port 9 nsew signal output
rlabel locali s 1516 333 1582 493 6 Y
port 9 nsew signal output
rlabel locali s 1348 333 1414 493 6 Y
port 9 nsew signal output
rlabel locali s 1012 333 1078 493 6 Y
port 9 nsew signal output
rlabel locali s 844 333 910 493 6 Y
port 9 nsew signal output
rlabel locali s 676 333 742 493 6 Y
port 9 nsew signal output
rlabel locali s 508 333 558 493 6 Y
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 2024 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1958780
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1943792
<< end >>
