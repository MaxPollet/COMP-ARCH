magic
tech sky130A
magscale 1 2
timestamp 1681267127
<< nwell >>
rect -38 261 590 582
<< pwell >>
rect 269 163 551 203
rect 4 27 551 163
rect 29 -17 63 27
rect 272 21 551 27
<< scnmos >>
rect 82 53 112 137
rect 154 53 184 137
rect 235 53 265 137
rect 356 47 386 177
rect 440 47 470 177
<< scpmoshvt >>
rect 81 311 111 395
rect 165 311 195 395
rect 260 297 290 381
rect 359 297 389 497
rect 443 297 473 497
<< ndiff >>
rect 295 137 356 177
rect 30 111 82 137
rect 30 77 38 111
rect 72 77 82 111
rect 30 53 82 77
rect 112 53 154 137
rect 184 53 235 137
rect 265 116 356 137
rect 265 82 311 116
rect 345 82 356 116
rect 265 53 356 82
rect 298 47 356 53
rect 386 123 440 177
rect 386 89 396 123
rect 430 89 440 123
rect 386 47 440 89
rect 470 120 525 177
rect 470 86 480 120
rect 514 86 525 120
rect 470 47 525 86
<< pdiff >>
rect 305 477 359 497
rect 305 443 315 477
rect 349 443 359 477
rect 305 408 359 443
rect 29 369 81 395
rect 29 335 37 369
rect 71 335 81 369
rect 29 311 81 335
rect 111 387 165 395
rect 111 353 121 387
rect 155 353 165 387
rect 111 311 165 353
rect 195 381 245 395
rect 305 381 315 408
rect 195 362 260 381
rect 195 328 216 362
rect 250 328 260 362
rect 195 311 260 328
rect 210 297 260 311
rect 290 374 315 381
rect 349 374 359 408
rect 290 297 359 374
rect 389 477 443 497
rect 389 443 399 477
rect 433 443 443 477
rect 389 409 443 443
rect 389 375 399 409
rect 433 375 443 409
rect 389 297 443 375
rect 473 477 525 497
rect 473 443 483 477
rect 517 443 525 477
rect 473 409 525 443
rect 473 375 483 409
rect 517 375 525 409
rect 473 297 525 375
<< ndiffc >>
rect 38 77 72 111
rect 311 82 345 116
rect 396 89 430 123
rect 480 86 514 120
<< pdiffc >>
rect 315 443 349 477
rect 37 335 71 369
rect 121 353 155 387
rect 216 328 250 362
rect 315 374 349 408
rect 399 443 433 477
rect 399 375 433 409
rect 483 443 517 477
rect 483 375 517 409
<< poly >>
rect 165 477 223 500
rect 165 443 179 477
rect 213 443 223 477
rect 165 427 223 443
rect 28 249 112 265
rect 28 215 38 249
rect 72 215 112 249
rect 28 199 112 215
rect 235 249 292 265
rect 235 215 245 249
rect 279 215 292 249
rect 235 199 292 215
rect 334 249 474 265
rect 334 215 344 249
rect 378 215 474 249
rect 334 199 474 215
<< polycont >>
rect 179 443 213 477
rect 38 215 72 249
rect 245 215 279 249
rect 344 215 378 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 17 426 143 527
rect 20 369 71 392
rect 20 335 37 369
rect 105 391 143 426
rect 179 477 274 493
rect 213 443 274 477
rect 179 425 274 443
rect 311 477 354 527
rect 311 443 315 477
rect 349 443 354 477
rect 311 408 354 443
rect 105 387 171 391
rect 105 353 121 387
rect 155 353 171 387
rect 216 362 266 378
rect 20 319 71 335
rect 250 328 266 362
rect 311 374 315 408
rect 349 374 354 408
rect 311 358 354 374
rect 394 477 449 493
rect 394 443 399 477
rect 433 443 449 477
rect 394 409 449 443
rect 394 375 399 409
rect 433 375 449 409
rect 394 359 449 375
rect 216 319 266 328
rect 20 285 378 319
rect 415 289 449 359
rect 483 477 535 527
rect 517 443 535 477
rect 483 409 535 443
rect 517 375 535 409
rect 483 325 535 375
rect 17 215 38 249
rect 72 215 94 249
rect 17 153 94 215
rect 128 114 179 285
rect 332 249 378 285
rect 21 111 179 114
rect 21 77 38 111
rect 72 77 179 111
rect 21 61 179 77
rect 213 215 245 249
rect 279 215 295 249
rect 213 150 295 215
rect 332 215 344 249
rect 332 199 378 215
rect 412 185 535 289
rect 213 61 259 150
rect 412 143 446 185
rect 396 123 446 143
rect 295 82 311 116
rect 345 82 361 116
rect 295 17 361 82
rect 430 89 446 123
rect 396 51 446 89
rect 480 120 535 149
rect 514 86 535 120
rect 480 17 535 86
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
<< metal1 >>
rect 0 561 552 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 0 496 552 527
rect 0 17 552 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
rect 0 -48 552 -17
<< labels >>
flabel locali s 213 425 247 459 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel locali s 397 85 431 119 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel locali s 397 425 431 459 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel locali s 29 153 63 187 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 213 153 247 187 0 FreeSans 400 0 0 0 C
port 3 nsew signal input
flabel locali s 489 221 523 255 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 46 544 46 544 0 FreeSans 200 0 0 0 VPWR
flabel metal1 s 46 0 46 0 0 FreeSans 200 0 0 0 VGND
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 and3_2
rlabel metal1 s 0 -48 552 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 552 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 552 544
string GDS_END 3858566
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3852742
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
