magic
tech sky130A
magscale 1 2
timestamp 1681267127
use sky130_fd_pr__hvdfm1sd__example_5595914180846  sky130_fd_pr__hvdfm1sd__example_5595914180846_0
timestamp 1681267127
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd__example_5595914180846  sky130_fd_pr__hvdfm1sd__example_5595914180846_1
timestamp 1681267127
transform 1 0 100 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 47708040
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 47706986
<< end >>
