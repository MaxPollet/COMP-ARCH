magic
tech sky130A
magscale 1 2
timestamp 1681267127
use sky130_fd_pr__dfm1sd__example_55959141808212  sky130_fd_pr__dfm1sd__example_55959141808212_0
timestamp 1681267127
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfm1sd__example_55959141808212  sky130_fd_pr__dfm1sd__example_55959141808212_1
timestamp 1681267127
transform 1 0 568 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_5595914180849  sky130_fd_pr__hvdfm1sd2__example_5595914180849_0
timestamp 1681267127
transform 1 0 100 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_5595914180849  sky130_fd_pr__hvdfm1sd2__example_5595914180849_1
timestamp 1681267127
transform 1 0 256 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_5595914180849  sky130_fd_pr__hvdfm1sd2__example_5595914180849_2
timestamp 1681267127
transform 1 0 412 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 37293740
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 37291142
<< end >>
