magic
tech sky130A
magscale 1 2
timestamp 1681267127
<< nwell >>
rect 726 -5168 1396 5168
<< pwell >>
rect 160 5320 1962 5766
rect 160 -5320 606 5320
rect 1516 -5320 1962 5320
rect 160 -5766 1962 -5320
<< mvpsubdiff >>
rect 186 5730 1936 5740
rect 186 5356 704 5730
rect 1418 5356 1936 5730
rect 186 5346 1936 5356
rect 186 5219 580 5346
rect 186 -5219 196 5219
rect 570 -5219 580 5219
rect 1542 5219 1936 5346
rect 186 -5346 580 -5219
rect 1542 -5219 1552 5219
rect 1926 -5219 1936 5219
rect 1542 -5346 1936 -5219
rect 186 -5356 1936 -5346
rect 186 -5730 704 -5356
rect 1418 -5730 1936 -5356
rect 186 -5740 1936 -5730
<< mvnsubdiff >>
rect 792 5068 945 5102
rect 979 5068 1013 5102
rect 1047 5068 1081 5102
rect 1115 5068 1149 5102
rect 1183 5068 1330 5102
rect 792 5015 896 5068
rect 792 4981 862 5015
rect 1232 5015 1330 5068
rect 792 4947 896 4981
rect 792 4913 862 4947
rect 792 4879 896 4913
rect 792 4845 862 4879
rect 792 4811 896 4845
rect 792 4777 862 4811
rect 792 4743 896 4777
rect 792 4709 862 4743
rect 792 4675 896 4709
rect 792 4641 862 4675
rect 792 4607 896 4641
rect 792 4573 862 4607
rect 792 4539 896 4573
rect 792 4505 862 4539
rect 792 4471 896 4505
rect 792 4437 862 4471
rect 792 4403 896 4437
rect 792 4369 862 4403
rect 792 4335 896 4369
rect 792 4301 862 4335
rect 792 4267 896 4301
rect 792 4233 862 4267
rect 792 4199 896 4233
rect 792 4165 862 4199
rect 792 4131 896 4165
rect 792 4097 862 4131
rect 792 4063 896 4097
rect 792 4029 862 4063
rect 792 3995 896 4029
rect 792 3961 862 3995
rect 792 3927 896 3961
rect 792 3893 862 3927
rect 792 3859 896 3893
rect 792 3825 862 3859
rect 792 3791 896 3825
rect 792 3757 862 3791
rect 792 3723 896 3757
rect 792 3689 862 3723
rect 792 3655 896 3689
rect 792 3621 862 3655
rect 792 3587 896 3621
rect 792 3553 862 3587
rect 792 3519 896 3553
rect 792 3485 862 3519
rect 792 3451 896 3485
rect 792 3417 862 3451
rect 792 3383 896 3417
rect 792 3349 862 3383
rect 792 3315 896 3349
rect 792 3281 862 3315
rect 792 3247 896 3281
rect 792 3213 862 3247
rect 792 3179 896 3213
rect 792 3145 862 3179
rect 792 3111 896 3145
rect 792 3077 862 3111
rect 792 3043 896 3077
rect 792 3009 862 3043
rect 792 2975 896 3009
rect 792 2941 862 2975
rect 792 2907 896 2941
rect 792 2873 862 2907
rect 792 2839 896 2873
rect 792 2805 862 2839
rect 792 2771 896 2805
rect 792 2737 862 2771
rect 792 2703 896 2737
rect 792 2669 862 2703
rect 792 2635 896 2669
rect 792 2601 862 2635
rect 792 2567 896 2601
rect 792 2533 862 2567
rect 792 2499 896 2533
rect 792 2465 862 2499
rect 792 2431 896 2465
rect 792 2397 862 2431
rect 792 2363 896 2397
rect 792 2329 862 2363
rect 792 2295 896 2329
rect 792 2261 862 2295
rect 792 2227 896 2261
rect 792 2193 862 2227
rect 792 2159 896 2193
rect 792 2125 862 2159
rect 792 2091 896 2125
rect 792 2057 862 2091
rect 792 2023 896 2057
rect 792 1989 862 2023
rect 792 1955 896 1989
rect 792 1921 862 1955
rect 792 1887 896 1921
rect 792 1853 862 1887
rect 792 1819 896 1853
rect 792 1785 862 1819
rect 792 1751 896 1785
rect 792 1717 862 1751
rect 792 1683 896 1717
rect 792 1649 862 1683
rect 792 1615 896 1649
rect 792 1581 862 1615
rect 792 1547 896 1581
rect 792 1513 862 1547
rect 792 1479 896 1513
rect 792 1445 862 1479
rect 792 1411 896 1445
rect 792 1377 862 1411
rect 792 1343 896 1377
rect 792 1309 862 1343
rect 792 1275 896 1309
rect 792 1241 862 1275
rect 792 1207 896 1241
rect 792 1173 862 1207
rect 792 1139 896 1173
rect 792 1105 862 1139
rect 792 1071 896 1105
rect 792 1037 862 1071
rect 792 1003 896 1037
rect 792 969 862 1003
rect 792 935 896 969
rect 792 901 862 935
rect 792 867 896 901
rect 792 833 862 867
rect 792 799 896 833
rect 792 765 862 799
rect 792 731 896 765
rect 792 697 862 731
rect 792 663 896 697
rect 792 629 862 663
rect 792 595 896 629
rect 792 561 862 595
rect 792 527 896 561
rect 792 493 862 527
rect 792 459 896 493
rect 792 425 862 459
rect 792 391 896 425
rect 792 357 862 391
rect 792 323 896 357
rect 792 289 862 323
rect 792 255 896 289
rect 792 221 862 255
rect 792 187 896 221
rect 792 153 862 187
rect 792 119 896 153
rect 792 85 862 119
rect 792 51 896 85
rect 792 17 862 51
rect 792 -17 896 17
rect 792 -51 862 -17
rect 792 -85 896 -51
rect 792 -119 862 -85
rect 792 -153 896 -119
rect 792 -187 862 -153
rect 792 -221 896 -187
rect 792 -255 862 -221
rect 792 -289 896 -255
rect 792 -323 862 -289
rect 792 -357 896 -323
rect 792 -391 862 -357
rect 792 -425 896 -391
rect 792 -459 862 -425
rect 792 -493 896 -459
rect 792 -527 862 -493
rect 792 -561 896 -527
rect 792 -595 862 -561
rect 792 -629 896 -595
rect 792 -663 862 -629
rect 792 -697 896 -663
rect 792 -731 862 -697
rect 792 -765 896 -731
rect 792 -799 862 -765
rect 792 -833 896 -799
rect 792 -867 862 -833
rect 792 -901 896 -867
rect 792 -935 862 -901
rect 792 -969 896 -935
rect 792 -1003 862 -969
rect 792 -1037 896 -1003
rect 792 -1071 862 -1037
rect 792 -1105 896 -1071
rect 792 -1139 862 -1105
rect 792 -1173 896 -1139
rect 792 -1207 862 -1173
rect 792 -1241 896 -1207
rect 792 -1275 862 -1241
rect 792 -1309 896 -1275
rect 792 -1343 862 -1309
rect 792 -1377 896 -1343
rect 792 -1411 862 -1377
rect 792 -1445 896 -1411
rect 792 -1479 862 -1445
rect 792 -1513 896 -1479
rect 792 -1547 862 -1513
rect 792 -1581 896 -1547
rect 792 -1615 862 -1581
rect 792 -1649 896 -1615
rect 792 -1683 862 -1649
rect 792 -1717 896 -1683
rect 792 -1751 862 -1717
rect 792 -1785 896 -1751
rect 792 -1819 862 -1785
rect 792 -1853 896 -1819
rect 792 -1887 862 -1853
rect 792 -1921 896 -1887
rect 792 -1955 862 -1921
rect 792 -1989 896 -1955
rect 792 -2023 862 -1989
rect 792 -2057 896 -2023
rect 792 -2091 862 -2057
rect 792 -2125 896 -2091
rect 792 -2159 862 -2125
rect 792 -2193 896 -2159
rect 792 -2227 862 -2193
rect 792 -2261 896 -2227
rect 792 -2295 862 -2261
rect 792 -2329 896 -2295
rect 792 -2363 862 -2329
rect 792 -2397 896 -2363
rect 792 -2431 862 -2397
rect 792 -2465 896 -2431
rect 792 -2499 862 -2465
rect 792 -2533 896 -2499
rect 792 -2567 862 -2533
rect 792 -2601 896 -2567
rect 792 -2635 862 -2601
rect 792 -2669 896 -2635
rect 792 -2703 862 -2669
rect 792 -2737 896 -2703
rect 792 -2771 862 -2737
rect 792 -2805 896 -2771
rect 792 -2839 862 -2805
rect 792 -2873 896 -2839
rect 792 -2907 862 -2873
rect 792 -2941 896 -2907
rect 792 -2975 862 -2941
rect 792 -3009 896 -2975
rect 792 -3043 862 -3009
rect 792 -3077 896 -3043
rect 792 -3111 862 -3077
rect 792 -3145 896 -3111
rect 792 -3179 862 -3145
rect 792 -3213 896 -3179
rect 792 -3247 862 -3213
rect 792 -3281 896 -3247
rect 792 -3315 862 -3281
rect 792 -3349 896 -3315
rect 792 -3383 862 -3349
rect 792 -3417 896 -3383
rect 792 -3451 862 -3417
rect 792 -3485 896 -3451
rect 792 -3519 862 -3485
rect 792 -3553 896 -3519
rect 792 -3587 862 -3553
rect 792 -3621 896 -3587
rect 792 -3655 862 -3621
rect 792 -3689 896 -3655
rect 792 -3723 862 -3689
rect 792 -3757 896 -3723
rect 792 -3791 862 -3757
rect 792 -3825 896 -3791
rect 792 -3859 862 -3825
rect 792 -3893 896 -3859
rect 792 -3927 862 -3893
rect 792 -3961 896 -3927
rect 792 -3995 862 -3961
rect 792 -4029 896 -3995
rect 792 -4063 862 -4029
rect 792 -4097 896 -4063
rect 792 -4131 862 -4097
rect 792 -4165 896 -4131
rect 792 -4199 862 -4165
rect 792 -4233 896 -4199
rect 792 -4267 862 -4233
rect 792 -4301 896 -4267
rect 792 -4335 862 -4301
rect 792 -4369 896 -4335
rect 792 -4403 862 -4369
rect 792 -4437 896 -4403
rect 792 -4471 862 -4437
rect 792 -4505 896 -4471
rect 792 -4539 862 -4505
rect 792 -4573 896 -4539
rect 792 -4607 862 -4573
rect 792 -4641 896 -4607
rect 792 -4675 862 -4641
rect 792 -4709 896 -4675
rect 792 -4743 862 -4709
rect 792 -4777 896 -4743
rect 792 -4811 862 -4777
rect 792 -4845 896 -4811
rect 792 -4879 862 -4845
rect 792 -4913 896 -4879
rect 792 -4947 862 -4913
rect 792 -4981 896 -4947
rect 792 -5015 862 -4981
rect 1266 4981 1330 5015
rect 1232 4947 1330 4981
rect 1266 4913 1330 4947
rect 1232 4879 1330 4913
rect 1266 4845 1330 4879
rect 1232 4811 1330 4845
rect 1266 4777 1330 4811
rect 1232 4743 1330 4777
rect 1266 4709 1330 4743
rect 1232 4675 1330 4709
rect 1266 4641 1330 4675
rect 1232 4607 1330 4641
rect 1266 4573 1330 4607
rect 1232 4539 1330 4573
rect 1266 4505 1330 4539
rect 1232 4471 1330 4505
rect 1266 4437 1330 4471
rect 1232 4403 1330 4437
rect 1266 4369 1330 4403
rect 1232 4335 1330 4369
rect 1266 4301 1330 4335
rect 1232 4267 1330 4301
rect 1266 4233 1330 4267
rect 1232 4199 1330 4233
rect 1266 4165 1330 4199
rect 1232 4131 1330 4165
rect 1266 4097 1330 4131
rect 1232 4063 1330 4097
rect 1266 4029 1330 4063
rect 1232 3995 1330 4029
rect 1266 3961 1330 3995
rect 1232 3927 1330 3961
rect 1266 3893 1330 3927
rect 1232 3859 1330 3893
rect 1266 3825 1330 3859
rect 1232 3791 1330 3825
rect 1266 3757 1330 3791
rect 1232 3723 1330 3757
rect 1266 3689 1330 3723
rect 1232 3655 1330 3689
rect 1266 3621 1330 3655
rect 1232 3587 1330 3621
rect 1266 3553 1330 3587
rect 1232 3519 1330 3553
rect 1266 3485 1330 3519
rect 1232 3451 1330 3485
rect 1266 3417 1330 3451
rect 1232 3383 1330 3417
rect 1266 3349 1330 3383
rect 1232 3315 1330 3349
rect 1266 3281 1330 3315
rect 1232 3247 1330 3281
rect 1266 3213 1330 3247
rect 1232 3179 1330 3213
rect 1266 3145 1330 3179
rect 1232 3111 1330 3145
rect 1266 3077 1330 3111
rect 1232 3043 1330 3077
rect 1266 3009 1330 3043
rect 1232 2975 1330 3009
rect 1266 2941 1330 2975
rect 1232 2907 1330 2941
rect 1266 2873 1330 2907
rect 1232 2839 1330 2873
rect 1266 2805 1330 2839
rect 1232 2771 1330 2805
rect 1266 2737 1330 2771
rect 1232 2703 1330 2737
rect 1266 2669 1330 2703
rect 1232 2635 1330 2669
rect 1266 2601 1330 2635
rect 1232 2567 1330 2601
rect 1266 2533 1330 2567
rect 1232 2499 1330 2533
rect 1266 2465 1330 2499
rect 1232 2431 1330 2465
rect 1266 2397 1330 2431
rect 1232 2363 1330 2397
rect 1266 2329 1330 2363
rect 1232 2295 1330 2329
rect 1266 2261 1330 2295
rect 1232 2227 1330 2261
rect 1266 2193 1330 2227
rect 1232 2159 1330 2193
rect 1266 2125 1330 2159
rect 1232 2091 1330 2125
rect 1266 2057 1330 2091
rect 1232 2023 1330 2057
rect 1266 1989 1330 2023
rect 1232 1955 1330 1989
rect 1266 1921 1330 1955
rect 1232 1887 1330 1921
rect 1266 1853 1330 1887
rect 1232 1819 1330 1853
rect 1266 1785 1330 1819
rect 1232 1751 1330 1785
rect 1266 1717 1330 1751
rect 1232 1683 1330 1717
rect 1266 1649 1330 1683
rect 1232 1615 1330 1649
rect 1266 1581 1330 1615
rect 1232 1547 1330 1581
rect 1266 1513 1330 1547
rect 1232 1479 1330 1513
rect 1266 1445 1330 1479
rect 1232 1411 1330 1445
rect 1266 1377 1330 1411
rect 1232 1343 1330 1377
rect 1266 1309 1330 1343
rect 1232 1275 1330 1309
rect 1266 1241 1330 1275
rect 1232 1207 1330 1241
rect 1266 1173 1330 1207
rect 1232 1139 1330 1173
rect 1266 1105 1330 1139
rect 1232 1071 1330 1105
rect 1266 1037 1330 1071
rect 1232 1003 1330 1037
rect 1266 969 1330 1003
rect 1232 935 1330 969
rect 1266 901 1330 935
rect 1232 867 1330 901
rect 1266 833 1330 867
rect 1232 799 1330 833
rect 1266 765 1330 799
rect 1232 731 1330 765
rect 1266 697 1330 731
rect 1232 663 1330 697
rect 1266 629 1330 663
rect 1232 595 1330 629
rect 1266 561 1330 595
rect 1232 527 1330 561
rect 1266 493 1330 527
rect 1232 459 1330 493
rect 1266 425 1330 459
rect 1232 391 1330 425
rect 1266 357 1330 391
rect 1232 323 1330 357
rect 1266 289 1330 323
rect 1232 255 1330 289
rect 1266 221 1330 255
rect 1232 187 1330 221
rect 1266 153 1330 187
rect 1232 119 1330 153
rect 1266 85 1330 119
rect 1232 51 1330 85
rect 1266 17 1330 51
rect 1232 -17 1330 17
rect 1266 -51 1330 -17
rect 1232 -85 1330 -51
rect 1266 -119 1330 -85
rect 1232 -153 1330 -119
rect 1266 -187 1330 -153
rect 1232 -221 1330 -187
rect 1266 -255 1330 -221
rect 1232 -289 1330 -255
rect 1266 -323 1330 -289
rect 1232 -357 1330 -323
rect 1266 -391 1330 -357
rect 1232 -425 1330 -391
rect 1266 -459 1330 -425
rect 1232 -493 1330 -459
rect 1266 -527 1330 -493
rect 1232 -561 1330 -527
rect 1266 -595 1330 -561
rect 1232 -629 1330 -595
rect 1266 -663 1330 -629
rect 1232 -697 1330 -663
rect 1266 -731 1330 -697
rect 1232 -765 1330 -731
rect 1266 -799 1330 -765
rect 1232 -833 1330 -799
rect 1266 -867 1330 -833
rect 1232 -901 1330 -867
rect 1266 -935 1330 -901
rect 1232 -969 1330 -935
rect 1266 -1003 1330 -969
rect 1232 -1037 1330 -1003
rect 1266 -1071 1330 -1037
rect 1232 -1105 1330 -1071
rect 1266 -1139 1330 -1105
rect 1232 -1173 1330 -1139
rect 1266 -1207 1330 -1173
rect 1232 -1241 1330 -1207
rect 1266 -1275 1330 -1241
rect 1232 -1309 1330 -1275
rect 1266 -1343 1330 -1309
rect 1232 -1377 1330 -1343
rect 1266 -1411 1330 -1377
rect 1232 -1445 1330 -1411
rect 1266 -1479 1330 -1445
rect 1232 -1513 1330 -1479
rect 1266 -1547 1330 -1513
rect 1232 -1581 1330 -1547
rect 1266 -1615 1330 -1581
rect 1232 -1649 1330 -1615
rect 1266 -1683 1330 -1649
rect 1232 -1717 1330 -1683
rect 1266 -1751 1330 -1717
rect 1232 -1785 1330 -1751
rect 1266 -1819 1330 -1785
rect 1232 -1853 1330 -1819
rect 1266 -1887 1330 -1853
rect 1232 -1921 1330 -1887
rect 1266 -1955 1330 -1921
rect 1232 -1989 1330 -1955
rect 1266 -2023 1330 -1989
rect 1232 -2057 1330 -2023
rect 1266 -2091 1330 -2057
rect 1232 -2125 1330 -2091
rect 1266 -2159 1330 -2125
rect 1232 -2193 1330 -2159
rect 1266 -2227 1330 -2193
rect 1232 -2261 1330 -2227
rect 1266 -2295 1330 -2261
rect 1232 -2329 1330 -2295
rect 1266 -2363 1330 -2329
rect 1232 -2397 1330 -2363
rect 1266 -2431 1330 -2397
rect 1232 -2465 1330 -2431
rect 1266 -2499 1330 -2465
rect 1232 -2533 1330 -2499
rect 1266 -2567 1330 -2533
rect 1232 -2601 1330 -2567
rect 1266 -2635 1330 -2601
rect 1232 -2669 1330 -2635
rect 1266 -2703 1330 -2669
rect 1232 -2737 1330 -2703
rect 1266 -2771 1330 -2737
rect 1232 -2805 1330 -2771
rect 1266 -2839 1330 -2805
rect 1232 -2873 1330 -2839
rect 1266 -2907 1330 -2873
rect 1232 -2941 1330 -2907
rect 1266 -2975 1330 -2941
rect 1232 -3009 1330 -2975
rect 1266 -3043 1330 -3009
rect 1232 -3077 1330 -3043
rect 1266 -3111 1330 -3077
rect 1232 -3145 1330 -3111
rect 1266 -3179 1330 -3145
rect 1232 -3213 1330 -3179
rect 1266 -3247 1330 -3213
rect 1232 -3281 1330 -3247
rect 1266 -3315 1330 -3281
rect 1232 -3349 1330 -3315
rect 1266 -3383 1330 -3349
rect 1232 -3417 1330 -3383
rect 1266 -3451 1330 -3417
rect 1232 -3485 1330 -3451
rect 1266 -3519 1330 -3485
rect 1232 -3553 1330 -3519
rect 1266 -3587 1330 -3553
rect 1232 -3621 1330 -3587
rect 1266 -3655 1330 -3621
rect 1232 -3689 1330 -3655
rect 1266 -3723 1330 -3689
rect 1232 -3757 1330 -3723
rect 1266 -3791 1330 -3757
rect 1232 -3825 1330 -3791
rect 1266 -3859 1330 -3825
rect 1232 -3893 1330 -3859
rect 1266 -3927 1330 -3893
rect 1232 -3961 1330 -3927
rect 1266 -3995 1330 -3961
rect 1232 -4029 1330 -3995
rect 1266 -4063 1330 -4029
rect 1232 -4097 1330 -4063
rect 1266 -4131 1330 -4097
rect 1232 -4165 1330 -4131
rect 1266 -4199 1330 -4165
rect 1232 -4233 1330 -4199
rect 1266 -4267 1330 -4233
rect 1232 -4301 1330 -4267
rect 1266 -4335 1330 -4301
rect 1232 -4369 1330 -4335
rect 1266 -4403 1330 -4369
rect 1232 -4437 1330 -4403
rect 1266 -4471 1330 -4437
rect 1232 -4505 1330 -4471
rect 1266 -4539 1330 -4505
rect 1232 -4573 1330 -4539
rect 1266 -4607 1330 -4573
rect 1232 -4641 1330 -4607
rect 1266 -4675 1330 -4641
rect 1232 -4709 1330 -4675
rect 1266 -4743 1330 -4709
rect 1232 -4777 1330 -4743
rect 1266 -4811 1330 -4777
rect 1232 -4845 1330 -4811
rect 1266 -4879 1330 -4845
rect 1232 -4913 1330 -4879
rect 1266 -4947 1330 -4913
rect 1232 -4981 1330 -4947
rect 792 -5068 896 -5015
rect 1266 -5015 1330 -4981
rect 1232 -5068 1330 -5015
rect 792 -5102 945 -5068
rect 979 -5102 1013 -5068
rect 1047 -5102 1081 -5068
rect 1115 -5102 1149 -5068
rect 1183 -5102 1330 -5068
<< mvpsubdiffcont >>
rect 704 5356 1418 5730
rect 196 -5219 570 5219
rect 1552 -5219 1926 5219
rect 704 -5730 1418 -5356
<< mvnsubdiffcont >>
rect 945 5068 979 5102
rect 1013 5068 1047 5102
rect 1081 5068 1115 5102
rect 1149 5068 1183 5102
rect 862 4981 896 5015
rect 862 4913 896 4947
rect 862 4845 896 4879
rect 862 4777 896 4811
rect 862 4709 896 4743
rect 862 4641 896 4675
rect 862 4573 896 4607
rect 862 4505 896 4539
rect 862 4437 896 4471
rect 862 4369 896 4403
rect 862 4301 896 4335
rect 862 4233 896 4267
rect 862 4165 896 4199
rect 862 4097 896 4131
rect 862 4029 896 4063
rect 862 3961 896 3995
rect 862 3893 896 3927
rect 862 3825 896 3859
rect 862 3757 896 3791
rect 862 3689 896 3723
rect 862 3621 896 3655
rect 862 3553 896 3587
rect 862 3485 896 3519
rect 862 3417 896 3451
rect 862 3349 896 3383
rect 862 3281 896 3315
rect 862 3213 896 3247
rect 862 3145 896 3179
rect 862 3077 896 3111
rect 862 3009 896 3043
rect 862 2941 896 2975
rect 862 2873 896 2907
rect 862 2805 896 2839
rect 862 2737 896 2771
rect 862 2669 896 2703
rect 862 2601 896 2635
rect 862 2533 896 2567
rect 862 2465 896 2499
rect 862 2397 896 2431
rect 862 2329 896 2363
rect 862 2261 896 2295
rect 862 2193 896 2227
rect 862 2125 896 2159
rect 862 2057 896 2091
rect 862 1989 896 2023
rect 862 1921 896 1955
rect 862 1853 896 1887
rect 862 1785 896 1819
rect 862 1717 896 1751
rect 862 1649 896 1683
rect 862 1581 896 1615
rect 862 1513 896 1547
rect 862 1445 896 1479
rect 862 1377 896 1411
rect 862 1309 896 1343
rect 862 1241 896 1275
rect 862 1173 896 1207
rect 862 1105 896 1139
rect 862 1037 896 1071
rect 862 969 896 1003
rect 862 901 896 935
rect 862 833 896 867
rect 862 765 896 799
rect 862 697 896 731
rect 862 629 896 663
rect 862 561 896 595
rect 862 493 896 527
rect 862 425 896 459
rect 862 357 896 391
rect 862 289 896 323
rect 862 221 896 255
rect 862 153 896 187
rect 862 85 896 119
rect 862 17 896 51
rect 862 -51 896 -17
rect 862 -119 896 -85
rect 862 -187 896 -153
rect 862 -255 896 -221
rect 862 -323 896 -289
rect 862 -391 896 -357
rect 862 -459 896 -425
rect 862 -527 896 -493
rect 862 -595 896 -561
rect 862 -663 896 -629
rect 862 -731 896 -697
rect 862 -799 896 -765
rect 862 -867 896 -833
rect 862 -935 896 -901
rect 862 -1003 896 -969
rect 862 -1071 896 -1037
rect 862 -1139 896 -1105
rect 862 -1207 896 -1173
rect 862 -1275 896 -1241
rect 862 -1343 896 -1309
rect 862 -1411 896 -1377
rect 862 -1479 896 -1445
rect 862 -1547 896 -1513
rect 862 -1615 896 -1581
rect 862 -1683 896 -1649
rect 862 -1751 896 -1717
rect 862 -1819 896 -1785
rect 862 -1887 896 -1853
rect 862 -1955 896 -1921
rect 862 -2023 896 -1989
rect 862 -2091 896 -2057
rect 862 -2159 896 -2125
rect 862 -2227 896 -2193
rect 862 -2295 896 -2261
rect 862 -2363 896 -2329
rect 862 -2431 896 -2397
rect 862 -2499 896 -2465
rect 862 -2567 896 -2533
rect 862 -2635 896 -2601
rect 862 -2703 896 -2669
rect 862 -2771 896 -2737
rect 862 -2839 896 -2805
rect 862 -2907 896 -2873
rect 862 -2975 896 -2941
rect 862 -3043 896 -3009
rect 862 -3111 896 -3077
rect 862 -3179 896 -3145
rect 862 -3247 896 -3213
rect 862 -3315 896 -3281
rect 862 -3383 896 -3349
rect 862 -3451 896 -3417
rect 862 -3519 896 -3485
rect 862 -3587 896 -3553
rect 862 -3655 896 -3621
rect 862 -3723 896 -3689
rect 862 -3791 896 -3757
rect 862 -3859 896 -3825
rect 862 -3927 896 -3893
rect 862 -3995 896 -3961
rect 862 -4063 896 -4029
rect 862 -4131 896 -4097
rect 862 -4199 896 -4165
rect 862 -4267 896 -4233
rect 862 -4335 896 -4301
rect 862 -4403 896 -4369
rect 862 -4471 896 -4437
rect 862 -4539 896 -4505
rect 862 -4607 896 -4573
rect 862 -4675 896 -4641
rect 862 -4743 896 -4709
rect 862 -4811 896 -4777
rect 862 -4879 896 -4845
rect 862 -4947 896 -4913
rect 862 -5015 896 -4981
rect 1232 4981 1266 5015
rect 1232 4913 1266 4947
rect 1232 4845 1266 4879
rect 1232 4777 1266 4811
rect 1232 4709 1266 4743
rect 1232 4641 1266 4675
rect 1232 4573 1266 4607
rect 1232 4505 1266 4539
rect 1232 4437 1266 4471
rect 1232 4369 1266 4403
rect 1232 4301 1266 4335
rect 1232 4233 1266 4267
rect 1232 4165 1266 4199
rect 1232 4097 1266 4131
rect 1232 4029 1266 4063
rect 1232 3961 1266 3995
rect 1232 3893 1266 3927
rect 1232 3825 1266 3859
rect 1232 3757 1266 3791
rect 1232 3689 1266 3723
rect 1232 3621 1266 3655
rect 1232 3553 1266 3587
rect 1232 3485 1266 3519
rect 1232 3417 1266 3451
rect 1232 3349 1266 3383
rect 1232 3281 1266 3315
rect 1232 3213 1266 3247
rect 1232 3145 1266 3179
rect 1232 3077 1266 3111
rect 1232 3009 1266 3043
rect 1232 2941 1266 2975
rect 1232 2873 1266 2907
rect 1232 2805 1266 2839
rect 1232 2737 1266 2771
rect 1232 2669 1266 2703
rect 1232 2601 1266 2635
rect 1232 2533 1266 2567
rect 1232 2465 1266 2499
rect 1232 2397 1266 2431
rect 1232 2329 1266 2363
rect 1232 2261 1266 2295
rect 1232 2193 1266 2227
rect 1232 2125 1266 2159
rect 1232 2057 1266 2091
rect 1232 1989 1266 2023
rect 1232 1921 1266 1955
rect 1232 1853 1266 1887
rect 1232 1785 1266 1819
rect 1232 1717 1266 1751
rect 1232 1649 1266 1683
rect 1232 1581 1266 1615
rect 1232 1513 1266 1547
rect 1232 1445 1266 1479
rect 1232 1377 1266 1411
rect 1232 1309 1266 1343
rect 1232 1241 1266 1275
rect 1232 1173 1266 1207
rect 1232 1105 1266 1139
rect 1232 1037 1266 1071
rect 1232 969 1266 1003
rect 1232 901 1266 935
rect 1232 833 1266 867
rect 1232 765 1266 799
rect 1232 697 1266 731
rect 1232 629 1266 663
rect 1232 561 1266 595
rect 1232 493 1266 527
rect 1232 425 1266 459
rect 1232 357 1266 391
rect 1232 289 1266 323
rect 1232 221 1266 255
rect 1232 153 1266 187
rect 1232 85 1266 119
rect 1232 17 1266 51
rect 1232 -51 1266 -17
rect 1232 -119 1266 -85
rect 1232 -187 1266 -153
rect 1232 -255 1266 -221
rect 1232 -323 1266 -289
rect 1232 -391 1266 -357
rect 1232 -459 1266 -425
rect 1232 -527 1266 -493
rect 1232 -595 1266 -561
rect 1232 -663 1266 -629
rect 1232 -731 1266 -697
rect 1232 -799 1266 -765
rect 1232 -867 1266 -833
rect 1232 -935 1266 -901
rect 1232 -1003 1266 -969
rect 1232 -1071 1266 -1037
rect 1232 -1139 1266 -1105
rect 1232 -1207 1266 -1173
rect 1232 -1275 1266 -1241
rect 1232 -1343 1266 -1309
rect 1232 -1411 1266 -1377
rect 1232 -1479 1266 -1445
rect 1232 -1547 1266 -1513
rect 1232 -1615 1266 -1581
rect 1232 -1683 1266 -1649
rect 1232 -1751 1266 -1717
rect 1232 -1819 1266 -1785
rect 1232 -1887 1266 -1853
rect 1232 -1955 1266 -1921
rect 1232 -2023 1266 -1989
rect 1232 -2091 1266 -2057
rect 1232 -2159 1266 -2125
rect 1232 -2227 1266 -2193
rect 1232 -2295 1266 -2261
rect 1232 -2363 1266 -2329
rect 1232 -2431 1266 -2397
rect 1232 -2499 1266 -2465
rect 1232 -2567 1266 -2533
rect 1232 -2635 1266 -2601
rect 1232 -2703 1266 -2669
rect 1232 -2771 1266 -2737
rect 1232 -2839 1266 -2805
rect 1232 -2907 1266 -2873
rect 1232 -2975 1266 -2941
rect 1232 -3043 1266 -3009
rect 1232 -3111 1266 -3077
rect 1232 -3179 1266 -3145
rect 1232 -3247 1266 -3213
rect 1232 -3315 1266 -3281
rect 1232 -3383 1266 -3349
rect 1232 -3451 1266 -3417
rect 1232 -3519 1266 -3485
rect 1232 -3587 1266 -3553
rect 1232 -3655 1266 -3621
rect 1232 -3723 1266 -3689
rect 1232 -3791 1266 -3757
rect 1232 -3859 1266 -3825
rect 1232 -3927 1266 -3893
rect 1232 -3995 1266 -3961
rect 1232 -4063 1266 -4029
rect 1232 -4131 1266 -4097
rect 1232 -4199 1266 -4165
rect 1232 -4267 1266 -4233
rect 1232 -4335 1266 -4301
rect 1232 -4403 1266 -4369
rect 1232 -4471 1266 -4437
rect 1232 -4539 1266 -4505
rect 1232 -4607 1266 -4573
rect 1232 -4675 1266 -4641
rect 1232 -4743 1266 -4709
rect 1232 -4811 1266 -4777
rect 1232 -4879 1266 -4845
rect 1232 -4947 1266 -4913
rect 1232 -5015 1266 -4981
rect 945 -5102 979 -5068
rect 1013 -5102 1047 -5068
rect 1081 -5102 1115 -5068
rect 1149 -5102 1183 -5068
<< mvpdiode >>
rect 964 4981 1164 5000
rect 964 -4981 979 4981
rect 1149 -4981 1164 4981
rect 964 -5000 1164 -4981
<< mvpdiodec >>
rect 979 -4981 1149 4981
<< locali >>
rect 186 5346 684 5740
rect 1438 5346 1936 5740
rect 186 5295 1936 5346
rect 186 5237 629 5295
rect 580 -5237 629 5237
rect 1488 5237 1936 5295
rect 792 5102 1330 5168
rect 792 5068 945 5102
rect 1009 5068 1013 5102
rect 1115 5068 1119 5102
rect 1183 5068 1330 5102
rect 792 5015 896 5068
rect 792 4951 862 5015
rect 1232 5015 1330 5068
rect 792 4947 896 4951
rect 792 4845 862 4947
rect 792 4841 896 4845
rect 792 4777 862 4841
rect 792 4769 896 4777
rect 792 4709 862 4769
rect 792 4697 896 4709
rect 792 4641 862 4697
rect 792 4625 896 4641
rect 792 4573 862 4625
rect 792 4553 896 4573
rect 792 4505 862 4553
rect 792 4481 896 4505
rect 792 4437 862 4481
rect 792 4409 896 4437
rect 792 4369 862 4409
rect 792 4337 896 4369
rect 792 4301 862 4337
rect 792 4267 896 4301
rect 792 4231 862 4267
rect 792 4199 896 4231
rect 792 4159 862 4199
rect 792 4131 896 4159
rect 792 4087 862 4131
rect 792 4063 896 4087
rect 792 4015 862 4063
rect 792 3995 896 4015
rect 792 3943 862 3995
rect 792 3927 896 3943
rect 792 3871 862 3927
rect 792 3859 896 3871
rect 792 3799 862 3859
rect 792 3791 896 3799
rect 792 3727 862 3791
rect 792 3723 896 3727
rect 792 3621 862 3723
rect 792 3617 896 3621
rect 792 3553 862 3617
rect 792 3545 896 3553
rect 792 3485 862 3545
rect 792 3473 896 3485
rect 792 3417 862 3473
rect 792 3401 896 3417
rect 792 3349 862 3401
rect 792 3329 896 3349
rect 792 3281 862 3329
rect 792 3257 896 3281
rect 792 3213 862 3257
rect 792 3185 896 3213
rect 792 3145 862 3185
rect 792 3113 896 3145
rect 792 3077 862 3113
rect 792 3043 896 3077
rect 792 3007 862 3043
rect 792 2975 896 3007
rect 792 2935 862 2975
rect 792 2907 896 2935
rect 792 2863 862 2907
rect 792 2839 896 2863
rect 792 2791 862 2839
rect 792 2771 896 2791
rect 792 2719 862 2771
rect 792 2703 896 2719
rect 792 2647 862 2703
rect 792 2635 896 2647
rect 792 2575 862 2635
rect 792 2567 896 2575
rect 792 2503 862 2567
rect 792 2499 896 2503
rect 792 2397 862 2499
rect 792 2393 896 2397
rect 792 2329 862 2393
rect 792 2321 896 2329
rect 792 2261 862 2321
rect 792 2249 896 2261
rect 792 2193 862 2249
rect 792 2177 896 2193
rect 792 2125 862 2177
rect 792 2105 896 2125
rect 792 2057 862 2105
rect 792 2033 896 2057
rect 792 1989 862 2033
rect 792 1961 896 1989
rect 792 1921 862 1961
rect 792 1889 896 1921
rect 792 1853 862 1889
rect 792 1819 896 1853
rect 792 1783 862 1819
rect 792 1751 896 1783
rect 792 1711 862 1751
rect 792 1683 896 1711
rect 792 1639 862 1683
rect 792 1615 896 1639
rect 792 1567 862 1615
rect 792 1547 896 1567
rect 792 1495 862 1547
rect 792 1479 896 1495
rect 792 1423 862 1479
rect 792 1411 896 1423
rect 792 1351 862 1411
rect 792 1343 896 1351
rect 792 1279 862 1343
rect 792 1275 896 1279
rect 792 1173 862 1275
rect 792 1169 896 1173
rect 792 1105 862 1169
rect 792 1097 896 1105
rect 792 1037 862 1097
rect 792 1025 896 1037
rect 792 969 862 1025
rect 792 953 896 969
rect 792 901 862 953
rect 792 881 896 901
rect 792 833 862 881
rect 792 809 896 833
rect 792 765 862 809
rect 792 737 896 765
rect 792 697 862 737
rect 792 665 896 697
rect 792 629 862 665
rect 792 595 896 629
rect 792 559 862 595
rect 792 527 896 559
rect 792 487 862 527
rect 792 459 896 487
rect 792 415 862 459
rect 792 391 896 415
rect 792 343 862 391
rect 792 323 896 343
rect 792 271 862 323
rect 792 255 896 271
rect 792 199 862 255
rect 792 187 896 199
rect 792 127 862 187
rect 792 119 896 127
rect 792 55 862 119
rect 792 51 896 55
rect 792 -51 862 51
rect 792 -55 896 -51
rect 792 -119 862 -55
rect 792 -127 896 -119
rect 792 -187 862 -127
rect 792 -199 896 -187
rect 792 -255 862 -199
rect 792 -271 896 -255
rect 792 -323 862 -271
rect 792 -343 896 -323
rect 792 -391 862 -343
rect 792 -415 896 -391
rect 792 -459 862 -415
rect 792 -487 896 -459
rect 792 -527 862 -487
rect 792 -559 896 -527
rect 792 -595 862 -559
rect 792 -629 896 -595
rect 792 -665 862 -629
rect 792 -697 896 -665
rect 792 -737 862 -697
rect 792 -765 896 -737
rect 792 -809 862 -765
rect 792 -833 896 -809
rect 792 -881 862 -833
rect 792 -901 896 -881
rect 792 -953 862 -901
rect 792 -969 896 -953
rect 792 -1025 862 -969
rect 792 -1037 896 -1025
rect 792 -1097 862 -1037
rect 792 -1105 896 -1097
rect 792 -1169 862 -1105
rect 792 -1173 896 -1169
rect 792 -1275 862 -1173
rect 792 -1279 896 -1275
rect 792 -1343 862 -1279
rect 792 -1351 896 -1343
rect 792 -1411 862 -1351
rect 792 -1423 896 -1411
rect 792 -1479 862 -1423
rect 792 -1495 896 -1479
rect 792 -1547 862 -1495
rect 792 -1567 896 -1547
rect 792 -1615 862 -1567
rect 792 -1639 896 -1615
rect 792 -1683 862 -1639
rect 792 -1711 896 -1683
rect 792 -1751 862 -1711
rect 792 -1783 896 -1751
rect 792 -1819 862 -1783
rect 792 -1853 896 -1819
rect 792 -1889 862 -1853
rect 792 -1921 896 -1889
rect 792 -1961 862 -1921
rect 792 -1989 896 -1961
rect 792 -2033 862 -1989
rect 792 -2057 896 -2033
rect 792 -2105 862 -2057
rect 792 -2125 896 -2105
rect 792 -2177 862 -2125
rect 792 -2193 896 -2177
rect 792 -2249 862 -2193
rect 792 -2261 896 -2249
rect 792 -2321 862 -2261
rect 792 -2329 896 -2321
rect 792 -2393 862 -2329
rect 792 -2397 896 -2393
rect 792 -2499 862 -2397
rect 792 -2503 896 -2499
rect 792 -2567 862 -2503
rect 792 -2575 896 -2567
rect 792 -2635 862 -2575
rect 792 -2647 896 -2635
rect 792 -2703 862 -2647
rect 792 -2719 896 -2703
rect 792 -2771 862 -2719
rect 792 -2791 896 -2771
rect 792 -2839 862 -2791
rect 792 -2863 896 -2839
rect 792 -2907 862 -2863
rect 792 -2935 896 -2907
rect 792 -2975 862 -2935
rect 792 -3007 896 -2975
rect 792 -3043 862 -3007
rect 792 -3077 896 -3043
rect 792 -3113 862 -3077
rect 792 -3145 896 -3113
rect 792 -3185 862 -3145
rect 792 -3213 896 -3185
rect 792 -3257 862 -3213
rect 792 -3281 896 -3257
rect 792 -3329 862 -3281
rect 792 -3349 896 -3329
rect 792 -3401 862 -3349
rect 792 -3417 896 -3401
rect 792 -3473 862 -3417
rect 792 -3485 896 -3473
rect 792 -3545 862 -3485
rect 792 -3553 896 -3545
rect 792 -3617 862 -3553
rect 792 -3621 896 -3617
rect 792 -3723 862 -3621
rect 792 -3727 896 -3723
rect 792 -3791 862 -3727
rect 792 -3799 896 -3791
rect 792 -3859 862 -3799
rect 792 -3871 896 -3859
rect 792 -3927 862 -3871
rect 792 -3943 896 -3927
rect 792 -3995 862 -3943
rect 792 -4015 896 -3995
rect 792 -4063 862 -4015
rect 792 -4087 896 -4063
rect 792 -4131 862 -4087
rect 792 -4159 896 -4131
rect 792 -4199 862 -4159
rect 792 -4231 896 -4199
rect 792 -4267 862 -4231
rect 792 -4301 896 -4267
rect 792 -4337 862 -4301
rect 792 -4369 896 -4337
rect 792 -4409 862 -4369
rect 792 -4437 896 -4409
rect 792 -4481 862 -4437
rect 792 -4505 896 -4481
rect 792 -4553 862 -4505
rect 792 -4573 896 -4553
rect 792 -4625 862 -4573
rect 792 -4641 896 -4625
rect 792 -4697 862 -4641
rect 792 -4709 896 -4697
rect 792 -4769 862 -4709
rect 792 -4777 896 -4769
rect 792 -4841 862 -4777
rect 792 -4845 896 -4841
rect 792 -4947 862 -4845
rect 792 -4951 896 -4947
rect 792 -5015 862 -4951
rect 976 4985 1152 5004
rect 976 4981 1011 4985
rect 1117 4981 1152 4985
rect 976 -4981 979 4981
rect 1149 -4981 1152 4981
rect 976 -4985 1011 -4981
rect 1117 -4985 1152 -4981
rect 976 -5004 1152 -4985
rect 1266 4951 1330 5015
rect 1232 4947 1330 4951
rect 1266 4845 1330 4947
rect 1232 4841 1330 4845
rect 1266 4777 1330 4841
rect 1232 4769 1330 4777
rect 1266 4709 1330 4769
rect 1232 4697 1330 4709
rect 1266 4641 1330 4697
rect 1232 4625 1330 4641
rect 1266 4573 1330 4625
rect 1232 4553 1330 4573
rect 1266 4505 1330 4553
rect 1232 4481 1330 4505
rect 1266 4437 1330 4481
rect 1232 4409 1330 4437
rect 1266 4369 1330 4409
rect 1232 4337 1330 4369
rect 1266 4301 1330 4337
rect 1232 4267 1330 4301
rect 1266 4231 1330 4267
rect 1232 4199 1330 4231
rect 1266 4159 1330 4199
rect 1232 4131 1330 4159
rect 1266 4087 1330 4131
rect 1232 4063 1330 4087
rect 1266 4015 1330 4063
rect 1232 3995 1330 4015
rect 1266 3943 1330 3995
rect 1232 3927 1330 3943
rect 1266 3871 1330 3927
rect 1232 3859 1330 3871
rect 1266 3799 1330 3859
rect 1232 3791 1330 3799
rect 1266 3727 1330 3791
rect 1232 3723 1330 3727
rect 1266 3621 1330 3723
rect 1232 3617 1330 3621
rect 1266 3553 1330 3617
rect 1232 3545 1330 3553
rect 1266 3485 1330 3545
rect 1232 3473 1330 3485
rect 1266 3417 1330 3473
rect 1232 3401 1330 3417
rect 1266 3349 1330 3401
rect 1232 3329 1330 3349
rect 1266 3281 1330 3329
rect 1232 3257 1330 3281
rect 1266 3213 1330 3257
rect 1232 3185 1330 3213
rect 1266 3145 1330 3185
rect 1232 3113 1330 3145
rect 1266 3077 1330 3113
rect 1232 3043 1330 3077
rect 1266 3007 1330 3043
rect 1232 2975 1330 3007
rect 1266 2935 1330 2975
rect 1232 2907 1330 2935
rect 1266 2863 1330 2907
rect 1232 2839 1330 2863
rect 1266 2791 1330 2839
rect 1232 2771 1330 2791
rect 1266 2719 1330 2771
rect 1232 2703 1330 2719
rect 1266 2647 1330 2703
rect 1232 2635 1330 2647
rect 1266 2575 1330 2635
rect 1232 2567 1330 2575
rect 1266 2503 1330 2567
rect 1232 2499 1330 2503
rect 1266 2397 1330 2499
rect 1232 2393 1330 2397
rect 1266 2329 1330 2393
rect 1232 2321 1330 2329
rect 1266 2261 1330 2321
rect 1232 2249 1330 2261
rect 1266 2193 1330 2249
rect 1232 2177 1330 2193
rect 1266 2125 1330 2177
rect 1232 2105 1330 2125
rect 1266 2057 1330 2105
rect 1232 2033 1330 2057
rect 1266 1989 1330 2033
rect 1232 1961 1330 1989
rect 1266 1921 1330 1961
rect 1232 1889 1330 1921
rect 1266 1853 1330 1889
rect 1232 1819 1330 1853
rect 1266 1783 1330 1819
rect 1232 1751 1330 1783
rect 1266 1711 1330 1751
rect 1232 1683 1330 1711
rect 1266 1639 1330 1683
rect 1232 1615 1330 1639
rect 1266 1567 1330 1615
rect 1232 1547 1330 1567
rect 1266 1495 1330 1547
rect 1232 1479 1330 1495
rect 1266 1423 1330 1479
rect 1232 1411 1330 1423
rect 1266 1351 1330 1411
rect 1232 1343 1330 1351
rect 1266 1279 1330 1343
rect 1232 1275 1330 1279
rect 1266 1173 1330 1275
rect 1232 1169 1330 1173
rect 1266 1105 1330 1169
rect 1232 1097 1330 1105
rect 1266 1037 1330 1097
rect 1232 1025 1330 1037
rect 1266 969 1330 1025
rect 1232 953 1330 969
rect 1266 901 1330 953
rect 1232 881 1330 901
rect 1266 833 1330 881
rect 1232 809 1330 833
rect 1266 765 1330 809
rect 1232 737 1330 765
rect 1266 697 1330 737
rect 1232 665 1330 697
rect 1266 629 1330 665
rect 1232 595 1330 629
rect 1266 559 1330 595
rect 1232 527 1330 559
rect 1266 487 1330 527
rect 1232 459 1330 487
rect 1266 415 1330 459
rect 1232 391 1330 415
rect 1266 343 1330 391
rect 1232 323 1330 343
rect 1266 271 1330 323
rect 1232 255 1330 271
rect 1266 199 1330 255
rect 1232 187 1330 199
rect 1266 127 1330 187
rect 1232 119 1330 127
rect 1266 55 1330 119
rect 1232 51 1330 55
rect 1266 -51 1330 51
rect 1232 -55 1330 -51
rect 1266 -119 1330 -55
rect 1232 -127 1330 -119
rect 1266 -187 1330 -127
rect 1232 -199 1330 -187
rect 1266 -255 1330 -199
rect 1232 -271 1330 -255
rect 1266 -323 1330 -271
rect 1232 -343 1330 -323
rect 1266 -391 1330 -343
rect 1232 -415 1330 -391
rect 1266 -459 1330 -415
rect 1232 -487 1330 -459
rect 1266 -527 1330 -487
rect 1232 -559 1330 -527
rect 1266 -595 1330 -559
rect 1232 -629 1330 -595
rect 1266 -665 1330 -629
rect 1232 -697 1330 -665
rect 1266 -737 1330 -697
rect 1232 -765 1330 -737
rect 1266 -809 1330 -765
rect 1232 -833 1330 -809
rect 1266 -881 1330 -833
rect 1232 -901 1330 -881
rect 1266 -953 1330 -901
rect 1232 -969 1330 -953
rect 1266 -1025 1330 -969
rect 1232 -1037 1330 -1025
rect 1266 -1097 1330 -1037
rect 1232 -1105 1330 -1097
rect 1266 -1169 1330 -1105
rect 1232 -1173 1330 -1169
rect 1266 -1275 1330 -1173
rect 1232 -1279 1330 -1275
rect 1266 -1343 1330 -1279
rect 1232 -1351 1330 -1343
rect 1266 -1411 1330 -1351
rect 1232 -1423 1330 -1411
rect 1266 -1479 1330 -1423
rect 1232 -1495 1330 -1479
rect 1266 -1547 1330 -1495
rect 1232 -1567 1330 -1547
rect 1266 -1615 1330 -1567
rect 1232 -1639 1330 -1615
rect 1266 -1683 1330 -1639
rect 1232 -1711 1330 -1683
rect 1266 -1751 1330 -1711
rect 1232 -1783 1330 -1751
rect 1266 -1819 1330 -1783
rect 1232 -1853 1330 -1819
rect 1266 -1889 1330 -1853
rect 1232 -1921 1330 -1889
rect 1266 -1961 1330 -1921
rect 1232 -1989 1330 -1961
rect 1266 -2033 1330 -1989
rect 1232 -2057 1330 -2033
rect 1266 -2105 1330 -2057
rect 1232 -2125 1330 -2105
rect 1266 -2177 1330 -2125
rect 1232 -2193 1330 -2177
rect 1266 -2249 1330 -2193
rect 1232 -2261 1330 -2249
rect 1266 -2321 1330 -2261
rect 1232 -2329 1330 -2321
rect 1266 -2393 1330 -2329
rect 1232 -2397 1330 -2393
rect 1266 -2499 1330 -2397
rect 1232 -2503 1330 -2499
rect 1266 -2567 1330 -2503
rect 1232 -2575 1330 -2567
rect 1266 -2635 1330 -2575
rect 1232 -2647 1330 -2635
rect 1266 -2703 1330 -2647
rect 1232 -2719 1330 -2703
rect 1266 -2771 1330 -2719
rect 1232 -2791 1330 -2771
rect 1266 -2839 1330 -2791
rect 1232 -2863 1330 -2839
rect 1266 -2907 1330 -2863
rect 1232 -2935 1330 -2907
rect 1266 -2975 1330 -2935
rect 1232 -3007 1330 -2975
rect 1266 -3043 1330 -3007
rect 1232 -3077 1330 -3043
rect 1266 -3113 1330 -3077
rect 1232 -3145 1330 -3113
rect 1266 -3185 1330 -3145
rect 1232 -3213 1330 -3185
rect 1266 -3257 1330 -3213
rect 1232 -3281 1330 -3257
rect 1266 -3329 1330 -3281
rect 1232 -3349 1330 -3329
rect 1266 -3401 1330 -3349
rect 1232 -3417 1330 -3401
rect 1266 -3473 1330 -3417
rect 1232 -3485 1330 -3473
rect 1266 -3545 1330 -3485
rect 1232 -3553 1330 -3545
rect 1266 -3617 1330 -3553
rect 1232 -3621 1330 -3617
rect 1266 -3723 1330 -3621
rect 1232 -3727 1330 -3723
rect 1266 -3791 1330 -3727
rect 1232 -3799 1330 -3791
rect 1266 -3859 1330 -3799
rect 1232 -3871 1330 -3859
rect 1266 -3927 1330 -3871
rect 1232 -3943 1330 -3927
rect 1266 -3995 1330 -3943
rect 1232 -4015 1330 -3995
rect 1266 -4063 1330 -4015
rect 1232 -4087 1330 -4063
rect 1266 -4131 1330 -4087
rect 1232 -4159 1330 -4131
rect 1266 -4199 1330 -4159
rect 1232 -4231 1330 -4199
rect 1266 -4267 1330 -4231
rect 1232 -4301 1330 -4267
rect 1266 -4337 1330 -4301
rect 1232 -4369 1330 -4337
rect 1266 -4409 1330 -4369
rect 1232 -4437 1330 -4409
rect 1266 -4481 1330 -4437
rect 1232 -4505 1330 -4481
rect 1266 -4553 1330 -4505
rect 1232 -4573 1330 -4553
rect 1266 -4625 1330 -4573
rect 1232 -4641 1330 -4625
rect 1266 -4697 1330 -4641
rect 1232 -4709 1330 -4697
rect 1266 -4769 1330 -4709
rect 1232 -4777 1330 -4769
rect 1266 -4841 1330 -4777
rect 1232 -4845 1330 -4841
rect 1266 -4947 1330 -4845
rect 1232 -4951 1330 -4947
rect 792 -5068 896 -5015
rect 1266 -5015 1330 -4951
rect 1232 -5068 1330 -5015
rect 792 -5102 945 -5068
rect 1009 -5102 1013 -5068
rect 1115 -5102 1119 -5068
rect 1183 -5102 1330 -5068
rect 792 -5168 1330 -5102
rect 186 -5286 629 -5237
rect 1488 -5237 1542 5237
rect 1488 -5286 1936 -5237
rect 186 -5346 1936 -5286
rect 186 -5740 684 -5346
rect 1438 -5740 1936 -5346
<< viali >>
rect 684 5730 1438 5740
rect 684 5356 704 5730
rect 704 5356 1418 5730
rect 1418 5356 1438 5730
rect 684 5346 1438 5356
rect 186 5219 580 5237
rect 186 -5219 196 5219
rect 196 -5219 570 5219
rect 570 -5219 580 5219
rect 186 -5237 580 -5219
rect 975 5068 979 5102
rect 979 5068 1009 5102
rect 1047 5068 1081 5102
rect 1119 5068 1149 5102
rect 1149 5068 1153 5102
rect 862 4981 896 4985
rect 862 4951 896 4981
rect 862 4879 896 4913
rect 862 4811 896 4841
rect 862 4807 896 4811
rect 862 4743 896 4769
rect 862 4735 896 4743
rect 862 4675 896 4697
rect 862 4663 896 4675
rect 862 4607 896 4625
rect 862 4591 896 4607
rect 862 4539 896 4553
rect 862 4519 896 4539
rect 862 4471 896 4481
rect 862 4447 896 4471
rect 862 4403 896 4409
rect 862 4375 896 4403
rect 862 4335 896 4337
rect 862 4303 896 4335
rect 862 4233 896 4265
rect 862 4231 896 4233
rect 862 4165 896 4193
rect 862 4159 896 4165
rect 862 4097 896 4121
rect 862 4087 896 4097
rect 862 4029 896 4049
rect 862 4015 896 4029
rect 862 3961 896 3977
rect 862 3943 896 3961
rect 862 3893 896 3905
rect 862 3871 896 3893
rect 862 3825 896 3833
rect 862 3799 896 3825
rect 862 3757 896 3761
rect 862 3727 896 3757
rect 862 3655 896 3689
rect 862 3587 896 3617
rect 862 3583 896 3587
rect 862 3519 896 3545
rect 862 3511 896 3519
rect 862 3451 896 3473
rect 862 3439 896 3451
rect 862 3383 896 3401
rect 862 3367 896 3383
rect 862 3315 896 3329
rect 862 3295 896 3315
rect 862 3247 896 3257
rect 862 3223 896 3247
rect 862 3179 896 3185
rect 862 3151 896 3179
rect 862 3111 896 3113
rect 862 3079 896 3111
rect 862 3009 896 3041
rect 862 3007 896 3009
rect 862 2941 896 2969
rect 862 2935 896 2941
rect 862 2873 896 2897
rect 862 2863 896 2873
rect 862 2805 896 2825
rect 862 2791 896 2805
rect 862 2737 896 2753
rect 862 2719 896 2737
rect 862 2669 896 2681
rect 862 2647 896 2669
rect 862 2601 896 2609
rect 862 2575 896 2601
rect 862 2533 896 2537
rect 862 2503 896 2533
rect 862 2431 896 2465
rect 862 2363 896 2393
rect 862 2359 896 2363
rect 862 2295 896 2321
rect 862 2287 896 2295
rect 862 2227 896 2249
rect 862 2215 896 2227
rect 862 2159 896 2177
rect 862 2143 896 2159
rect 862 2091 896 2105
rect 862 2071 896 2091
rect 862 2023 896 2033
rect 862 1999 896 2023
rect 862 1955 896 1961
rect 862 1927 896 1955
rect 862 1887 896 1889
rect 862 1855 896 1887
rect 862 1785 896 1817
rect 862 1783 896 1785
rect 862 1717 896 1745
rect 862 1711 896 1717
rect 862 1649 896 1673
rect 862 1639 896 1649
rect 862 1581 896 1601
rect 862 1567 896 1581
rect 862 1513 896 1529
rect 862 1495 896 1513
rect 862 1445 896 1457
rect 862 1423 896 1445
rect 862 1377 896 1385
rect 862 1351 896 1377
rect 862 1309 896 1313
rect 862 1279 896 1309
rect 862 1207 896 1241
rect 862 1139 896 1169
rect 862 1135 896 1139
rect 862 1071 896 1097
rect 862 1063 896 1071
rect 862 1003 896 1025
rect 862 991 896 1003
rect 862 935 896 953
rect 862 919 896 935
rect 862 867 896 881
rect 862 847 896 867
rect 862 799 896 809
rect 862 775 896 799
rect 862 731 896 737
rect 862 703 896 731
rect 862 663 896 665
rect 862 631 896 663
rect 862 561 896 593
rect 862 559 896 561
rect 862 493 896 521
rect 862 487 896 493
rect 862 425 896 449
rect 862 415 896 425
rect 862 357 896 377
rect 862 343 896 357
rect 862 289 896 305
rect 862 271 896 289
rect 862 221 896 233
rect 862 199 896 221
rect 862 153 896 161
rect 862 127 896 153
rect 862 85 896 89
rect 862 55 896 85
rect 862 -17 896 17
rect 862 -85 896 -55
rect 862 -89 896 -85
rect 862 -153 896 -127
rect 862 -161 896 -153
rect 862 -221 896 -199
rect 862 -233 896 -221
rect 862 -289 896 -271
rect 862 -305 896 -289
rect 862 -357 896 -343
rect 862 -377 896 -357
rect 862 -425 896 -415
rect 862 -449 896 -425
rect 862 -493 896 -487
rect 862 -521 896 -493
rect 862 -561 896 -559
rect 862 -593 896 -561
rect 862 -663 896 -631
rect 862 -665 896 -663
rect 862 -731 896 -703
rect 862 -737 896 -731
rect 862 -799 896 -775
rect 862 -809 896 -799
rect 862 -867 896 -847
rect 862 -881 896 -867
rect 862 -935 896 -919
rect 862 -953 896 -935
rect 862 -1003 896 -991
rect 862 -1025 896 -1003
rect 862 -1071 896 -1063
rect 862 -1097 896 -1071
rect 862 -1139 896 -1135
rect 862 -1169 896 -1139
rect 862 -1241 896 -1207
rect 862 -1309 896 -1279
rect 862 -1313 896 -1309
rect 862 -1377 896 -1351
rect 862 -1385 896 -1377
rect 862 -1445 896 -1423
rect 862 -1457 896 -1445
rect 862 -1513 896 -1495
rect 862 -1529 896 -1513
rect 862 -1581 896 -1567
rect 862 -1601 896 -1581
rect 862 -1649 896 -1639
rect 862 -1673 896 -1649
rect 862 -1717 896 -1711
rect 862 -1745 896 -1717
rect 862 -1785 896 -1783
rect 862 -1817 896 -1785
rect 862 -1887 896 -1855
rect 862 -1889 896 -1887
rect 862 -1955 896 -1927
rect 862 -1961 896 -1955
rect 862 -2023 896 -1999
rect 862 -2033 896 -2023
rect 862 -2091 896 -2071
rect 862 -2105 896 -2091
rect 862 -2159 896 -2143
rect 862 -2177 896 -2159
rect 862 -2227 896 -2215
rect 862 -2249 896 -2227
rect 862 -2295 896 -2287
rect 862 -2321 896 -2295
rect 862 -2363 896 -2359
rect 862 -2393 896 -2363
rect 862 -2465 896 -2431
rect 862 -2533 896 -2503
rect 862 -2537 896 -2533
rect 862 -2601 896 -2575
rect 862 -2609 896 -2601
rect 862 -2669 896 -2647
rect 862 -2681 896 -2669
rect 862 -2737 896 -2719
rect 862 -2753 896 -2737
rect 862 -2805 896 -2791
rect 862 -2825 896 -2805
rect 862 -2873 896 -2863
rect 862 -2897 896 -2873
rect 862 -2941 896 -2935
rect 862 -2969 896 -2941
rect 862 -3009 896 -3007
rect 862 -3041 896 -3009
rect 862 -3111 896 -3079
rect 862 -3113 896 -3111
rect 862 -3179 896 -3151
rect 862 -3185 896 -3179
rect 862 -3247 896 -3223
rect 862 -3257 896 -3247
rect 862 -3315 896 -3295
rect 862 -3329 896 -3315
rect 862 -3383 896 -3367
rect 862 -3401 896 -3383
rect 862 -3451 896 -3439
rect 862 -3473 896 -3451
rect 862 -3519 896 -3511
rect 862 -3545 896 -3519
rect 862 -3587 896 -3583
rect 862 -3617 896 -3587
rect 862 -3689 896 -3655
rect 862 -3757 896 -3727
rect 862 -3761 896 -3757
rect 862 -3825 896 -3799
rect 862 -3833 896 -3825
rect 862 -3893 896 -3871
rect 862 -3905 896 -3893
rect 862 -3961 896 -3943
rect 862 -3977 896 -3961
rect 862 -4029 896 -4015
rect 862 -4049 896 -4029
rect 862 -4097 896 -4087
rect 862 -4121 896 -4097
rect 862 -4165 896 -4159
rect 862 -4193 896 -4165
rect 862 -4233 896 -4231
rect 862 -4265 896 -4233
rect 862 -4335 896 -4303
rect 862 -4337 896 -4335
rect 862 -4403 896 -4375
rect 862 -4409 896 -4403
rect 862 -4471 896 -4447
rect 862 -4481 896 -4471
rect 862 -4539 896 -4519
rect 862 -4553 896 -4539
rect 862 -4607 896 -4591
rect 862 -4625 896 -4607
rect 862 -4675 896 -4663
rect 862 -4697 896 -4675
rect 862 -4743 896 -4735
rect 862 -4769 896 -4743
rect 862 -4811 896 -4807
rect 862 -4841 896 -4811
rect 862 -4913 896 -4879
rect 862 -4981 896 -4951
rect 862 -4985 896 -4981
rect 1011 4981 1117 4985
rect 1011 -4981 1117 4981
rect 1011 -4985 1117 -4981
rect 1232 4981 1266 4985
rect 1232 4951 1266 4981
rect 1232 4879 1266 4913
rect 1232 4811 1266 4841
rect 1232 4807 1266 4811
rect 1232 4743 1266 4769
rect 1232 4735 1266 4743
rect 1232 4675 1266 4697
rect 1232 4663 1266 4675
rect 1232 4607 1266 4625
rect 1232 4591 1266 4607
rect 1232 4539 1266 4553
rect 1232 4519 1266 4539
rect 1232 4471 1266 4481
rect 1232 4447 1266 4471
rect 1232 4403 1266 4409
rect 1232 4375 1266 4403
rect 1232 4335 1266 4337
rect 1232 4303 1266 4335
rect 1232 4233 1266 4265
rect 1232 4231 1266 4233
rect 1232 4165 1266 4193
rect 1232 4159 1266 4165
rect 1232 4097 1266 4121
rect 1232 4087 1266 4097
rect 1232 4029 1266 4049
rect 1232 4015 1266 4029
rect 1232 3961 1266 3977
rect 1232 3943 1266 3961
rect 1232 3893 1266 3905
rect 1232 3871 1266 3893
rect 1232 3825 1266 3833
rect 1232 3799 1266 3825
rect 1232 3757 1266 3761
rect 1232 3727 1266 3757
rect 1232 3655 1266 3689
rect 1232 3587 1266 3617
rect 1232 3583 1266 3587
rect 1232 3519 1266 3545
rect 1232 3511 1266 3519
rect 1232 3451 1266 3473
rect 1232 3439 1266 3451
rect 1232 3383 1266 3401
rect 1232 3367 1266 3383
rect 1232 3315 1266 3329
rect 1232 3295 1266 3315
rect 1232 3247 1266 3257
rect 1232 3223 1266 3247
rect 1232 3179 1266 3185
rect 1232 3151 1266 3179
rect 1232 3111 1266 3113
rect 1232 3079 1266 3111
rect 1232 3009 1266 3041
rect 1232 3007 1266 3009
rect 1232 2941 1266 2969
rect 1232 2935 1266 2941
rect 1232 2873 1266 2897
rect 1232 2863 1266 2873
rect 1232 2805 1266 2825
rect 1232 2791 1266 2805
rect 1232 2737 1266 2753
rect 1232 2719 1266 2737
rect 1232 2669 1266 2681
rect 1232 2647 1266 2669
rect 1232 2601 1266 2609
rect 1232 2575 1266 2601
rect 1232 2533 1266 2537
rect 1232 2503 1266 2533
rect 1232 2431 1266 2465
rect 1232 2363 1266 2393
rect 1232 2359 1266 2363
rect 1232 2295 1266 2321
rect 1232 2287 1266 2295
rect 1232 2227 1266 2249
rect 1232 2215 1266 2227
rect 1232 2159 1266 2177
rect 1232 2143 1266 2159
rect 1232 2091 1266 2105
rect 1232 2071 1266 2091
rect 1232 2023 1266 2033
rect 1232 1999 1266 2023
rect 1232 1955 1266 1961
rect 1232 1927 1266 1955
rect 1232 1887 1266 1889
rect 1232 1855 1266 1887
rect 1232 1785 1266 1817
rect 1232 1783 1266 1785
rect 1232 1717 1266 1745
rect 1232 1711 1266 1717
rect 1232 1649 1266 1673
rect 1232 1639 1266 1649
rect 1232 1581 1266 1601
rect 1232 1567 1266 1581
rect 1232 1513 1266 1529
rect 1232 1495 1266 1513
rect 1232 1445 1266 1457
rect 1232 1423 1266 1445
rect 1232 1377 1266 1385
rect 1232 1351 1266 1377
rect 1232 1309 1266 1313
rect 1232 1279 1266 1309
rect 1232 1207 1266 1241
rect 1232 1139 1266 1169
rect 1232 1135 1266 1139
rect 1232 1071 1266 1097
rect 1232 1063 1266 1071
rect 1232 1003 1266 1025
rect 1232 991 1266 1003
rect 1232 935 1266 953
rect 1232 919 1266 935
rect 1232 867 1266 881
rect 1232 847 1266 867
rect 1232 799 1266 809
rect 1232 775 1266 799
rect 1232 731 1266 737
rect 1232 703 1266 731
rect 1232 663 1266 665
rect 1232 631 1266 663
rect 1232 561 1266 593
rect 1232 559 1266 561
rect 1232 493 1266 521
rect 1232 487 1266 493
rect 1232 425 1266 449
rect 1232 415 1266 425
rect 1232 357 1266 377
rect 1232 343 1266 357
rect 1232 289 1266 305
rect 1232 271 1266 289
rect 1232 221 1266 233
rect 1232 199 1266 221
rect 1232 153 1266 161
rect 1232 127 1266 153
rect 1232 85 1266 89
rect 1232 55 1266 85
rect 1232 -17 1266 17
rect 1232 -85 1266 -55
rect 1232 -89 1266 -85
rect 1232 -153 1266 -127
rect 1232 -161 1266 -153
rect 1232 -221 1266 -199
rect 1232 -233 1266 -221
rect 1232 -289 1266 -271
rect 1232 -305 1266 -289
rect 1232 -357 1266 -343
rect 1232 -377 1266 -357
rect 1232 -425 1266 -415
rect 1232 -449 1266 -425
rect 1232 -493 1266 -487
rect 1232 -521 1266 -493
rect 1232 -561 1266 -559
rect 1232 -593 1266 -561
rect 1232 -663 1266 -631
rect 1232 -665 1266 -663
rect 1232 -731 1266 -703
rect 1232 -737 1266 -731
rect 1232 -799 1266 -775
rect 1232 -809 1266 -799
rect 1232 -867 1266 -847
rect 1232 -881 1266 -867
rect 1232 -935 1266 -919
rect 1232 -953 1266 -935
rect 1232 -1003 1266 -991
rect 1232 -1025 1266 -1003
rect 1232 -1071 1266 -1063
rect 1232 -1097 1266 -1071
rect 1232 -1139 1266 -1135
rect 1232 -1169 1266 -1139
rect 1232 -1241 1266 -1207
rect 1232 -1309 1266 -1279
rect 1232 -1313 1266 -1309
rect 1232 -1377 1266 -1351
rect 1232 -1385 1266 -1377
rect 1232 -1445 1266 -1423
rect 1232 -1457 1266 -1445
rect 1232 -1513 1266 -1495
rect 1232 -1529 1266 -1513
rect 1232 -1581 1266 -1567
rect 1232 -1601 1266 -1581
rect 1232 -1649 1266 -1639
rect 1232 -1673 1266 -1649
rect 1232 -1717 1266 -1711
rect 1232 -1745 1266 -1717
rect 1232 -1785 1266 -1783
rect 1232 -1817 1266 -1785
rect 1232 -1887 1266 -1855
rect 1232 -1889 1266 -1887
rect 1232 -1955 1266 -1927
rect 1232 -1961 1266 -1955
rect 1232 -2023 1266 -1999
rect 1232 -2033 1266 -2023
rect 1232 -2091 1266 -2071
rect 1232 -2105 1266 -2091
rect 1232 -2159 1266 -2143
rect 1232 -2177 1266 -2159
rect 1232 -2227 1266 -2215
rect 1232 -2249 1266 -2227
rect 1232 -2295 1266 -2287
rect 1232 -2321 1266 -2295
rect 1232 -2363 1266 -2359
rect 1232 -2393 1266 -2363
rect 1232 -2465 1266 -2431
rect 1232 -2533 1266 -2503
rect 1232 -2537 1266 -2533
rect 1232 -2601 1266 -2575
rect 1232 -2609 1266 -2601
rect 1232 -2669 1266 -2647
rect 1232 -2681 1266 -2669
rect 1232 -2737 1266 -2719
rect 1232 -2753 1266 -2737
rect 1232 -2805 1266 -2791
rect 1232 -2825 1266 -2805
rect 1232 -2873 1266 -2863
rect 1232 -2897 1266 -2873
rect 1232 -2941 1266 -2935
rect 1232 -2969 1266 -2941
rect 1232 -3009 1266 -3007
rect 1232 -3041 1266 -3009
rect 1232 -3111 1266 -3079
rect 1232 -3113 1266 -3111
rect 1232 -3179 1266 -3151
rect 1232 -3185 1266 -3179
rect 1232 -3247 1266 -3223
rect 1232 -3257 1266 -3247
rect 1232 -3315 1266 -3295
rect 1232 -3329 1266 -3315
rect 1232 -3383 1266 -3367
rect 1232 -3401 1266 -3383
rect 1232 -3451 1266 -3439
rect 1232 -3473 1266 -3451
rect 1232 -3519 1266 -3511
rect 1232 -3545 1266 -3519
rect 1232 -3587 1266 -3583
rect 1232 -3617 1266 -3587
rect 1232 -3689 1266 -3655
rect 1232 -3757 1266 -3727
rect 1232 -3761 1266 -3757
rect 1232 -3825 1266 -3799
rect 1232 -3833 1266 -3825
rect 1232 -3893 1266 -3871
rect 1232 -3905 1266 -3893
rect 1232 -3961 1266 -3943
rect 1232 -3977 1266 -3961
rect 1232 -4029 1266 -4015
rect 1232 -4049 1266 -4029
rect 1232 -4097 1266 -4087
rect 1232 -4121 1266 -4097
rect 1232 -4165 1266 -4159
rect 1232 -4193 1266 -4165
rect 1232 -4233 1266 -4231
rect 1232 -4265 1266 -4233
rect 1232 -4335 1266 -4303
rect 1232 -4337 1266 -4335
rect 1232 -4403 1266 -4375
rect 1232 -4409 1266 -4403
rect 1232 -4471 1266 -4447
rect 1232 -4481 1266 -4471
rect 1232 -4539 1266 -4519
rect 1232 -4553 1266 -4539
rect 1232 -4607 1266 -4591
rect 1232 -4625 1266 -4607
rect 1232 -4675 1266 -4663
rect 1232 -4697 1266 -4675
rect 1232 -4743 1266 -4735
rect 1232 -4769 1266 -4743
rect 1232 -4811 1266 -4807
rect 1232 -4841 1266 -4811
rect 1232 -4913 1266 -4879
rect 1232 -4981 1266 -4951
rect 1232 -4985 1266 -4981
rect 975 -5102 979 -5068
rect 979 -5102 1009 -5068
rect 1047 -5102 1081 -5068
rect 1119 -5102 1149 -5068
rect 1149 -5102 1153 -5068
rect 1542 5219 1936 5237
rect 1542 -5219 1552 5219
rect 1552 -5219 1926 5219
rect 1926 -5219 1936 5219
rect 1542 -5237 1936 -5219
rect 684 -5356 1438 -5346
rect 684 -5730 704 -5356
rect 704 -5730 1418 -5356
rect 1418 -5730 1438 -5356
rect 684 -5740 1438 -5730
<< metal1 >>
tri 546 5740 566 5760 se
rect 566 5740 1556 5760
tri 166 5360 546 5740 se
rect 546 5360 684 5740
rect 166 5346 684 5360
rect 1438 5360 1556 5740
tri 1556 5360 1956 5760 sw
rect 1438 5346 1956 5360
rect 166 5295 1956 5346
rect 166 5268 642 5295
tri 642 5268 669 5295 nw
tri 1448 5268 1475 5295 ne
rect 1475 5268 1956 5295
rect 166 5237 629 5268
tri 629 5255 642 5268 nw
tri 1475 5255 1488 5268 ne
rect 166 -5237 186 5237
rect 580 -5237 629 5237
rect 1488 5237 1956 5268
rect 792 5102 1330 5168
rect 792 5068 975 5102
rect 1009 5068 1047 5102
rect 1081 5068 1119 5102
rect 1153 5068 1330 5102
rect 792 5062 1330 5068
rect 792 4985 902 5062
tri 902 5022 942 5062 nw
tri 1186 5022 1226 5062 ne
rect 792 4951 862 4985
rect 896 4951 902 4985
rect 792 4913 902 4951
rect 792 4879 862 4913
rect 896 4879 902 4913
rect 792 4841 902 4879
rect 792 4807 862 4841
rect 896 4807 902 4841
rect 792 4769 902 4807
rect 792 4735 862 4769
rect 896 4735 902 4769
rect 792 4697 902 4735
rect 792 4663 862 4697
rect 896 4663 902 4697
rect 792 4625 902 4663
rect 792 4591 862 4625
rect 896 4591 902 4625
rect 792 4553 902 4591
rect 792 4519 862 4553
rect 896 4519 902 4553
rect 792 4481 902 4519
rect 792 4447 862 4481
rect 896 4447 902 4481
rect 792 4409 902 4447
rect 792 4375 862 4409
rect 896 4375 902 4409
rect 792 4337 902 4375
rect 792 4303 862 4337
rect 896 4303 902 4337
rect 792 4265 902 4303
rect 792 4231 862 4265
rect 896 4231 902 4265
rect 792 4193 902 4231
rect 792 4159 862 4193
rect 896 4159 902 4193
rect 792 4121 902 4159
rect 792 4087 862 4121
rect 896 4087 902 4121
rect 792 4049 902 4087
rect 792 4015 862 4049
rect 896 4015 902 4049
rect 792 3977 902 4015
rect 792 3943 862 3977
rect 896 3943 902 3977
rect 792 3905 902 3943
rect 792 3871 862 3905
rect 896 3871 902 3905
rect 792 3833 902 3871
rect 792 3799 862 3833
rect 896 3799 902 3833
rect 792 3761 902 3799
rect 792 3727 862 3761
rect 896 3727 902 3761
rect 792 3689 902 3727
rect 792 3655 862 3689
rect 896 3655 902 3689
rect 792 3617 902 3655
rect 792 3583 862 3617
rect 896 3583 902 3617
rect 792 3545 902 3583
rect 792 3511 862 3545
rect 896 3511 902 3545
rect 792 3473 902 3511
rect 792 3439 862 3473
rect 896 3439 902 3473
rect 792 3401 902 3439
rect 792 3367 862 3401
rect 896 3367 902 3401
rect 792 3329 902 3367
rect 792 3295 862 3329
rect 896 3295 902 3329
rect 792 3257 902 3295
rect 792 3223 862 3257
rect 896 3223 902 3257
rect 792 3185 902 3223
rect 792 3151 862 3185
rect 896 3151 902 3185
rect 792 3113 902 3151
rect 792 3079 862 3113
rect 896 3079 902 3113
rect 792 3041 902 3079
rect 792 3007 862 3041
rect 896 3007 902 3041
rect 792 2969 902 3007
rect 792 2935 862 2969
rect 896 2935 902 2969
rect 792 2897 902 2935
rect 792 2863 862 2897
rect 896 2863 902 2897
rect 792 2825 902 2863
rect 792 2791 862 2825
rect 896 2791 902 2825
rect 792 2753 902 2791
rect 792 2719 862 2753
rect 896 2719 902 2753
rect 792 2681 902 2719
rect 792 2647 862 2681
rect 896 2647 902 2681
rect 792 2609 902 2647
rect 792 2575 862 2609
rect 896 2575 902 2609
rect 792 2537 902 2575
rect 792 2503 862 2537
rect 896 2503 902 2537
rect 792 2465 902 2503
rect 792 2431 862 2465
rect 896 2431 902 2465
rect 792 2393 902 2431
rect 792 2359 862 2393
rect 896 2359 902 2393
rect 792 2321 902 2359
rect 792 2287 862 2321
rect 896 2287 902 2321
rect 792 2249 902 2287
rect 792 2215 862 2249
rect 896 2215 902 2249
rect 792 2177 902 2215
rect 792 2143 862 2177
rect 896 2143 902 2177
rect 792 2105 902 2143
rect 792 2071 862 2105
rect 896 2071 902 2105
rect 792 2033 902 2071
rect 792 1999 862 2033
rect 896 1999 902 2033
rect 792 1961 902 1999
rect 792 1927 862 1961
rect 896 1927 902 1961
rect 792 1889 902 1927
rect 792 1855 862 1889
rect 896 1855 902 1889
rect 792 1817 902 1855
rect 792 1783 862 1817
rect 896 1783 902 1817
rect 792 1745 902 1783
rect 792 1711 862 1745
rect 896 1711 902 1745
rect 792 1673 902 1711
rect 792 1639 862 1673
rect 896 1639 902 1673
rect 792 1601 902 1639
rect 792 1567 862 1601
rect 896 1567 902 1601
rect 792 1529 902 1567
rect 792 1495 862 1529
rect 896 1495 902 1529
rect 792 1457 902 1495
rect 792 1423 862 1457
rect 896 1423 902 1457
rect 792 1385 902 1423
rect 792 1351 862 1385
rect 896 1351 902 1385
rect 792 1313 902 1351
rect 792 1279 862 1313
rect 896 1279 902 1313
rect 792 1241 902 1279
rect 792 1207 862 1241
rect 896 1207 902 1241
rect 792 1169 902 1207
rect 792 1135 862 1169
rect 896 1135 902 1169
rect 792 1097 902 1135
rect 792 1063 862 1097
rect 896 1063 902 1097
rect 792 1025 902 1063
rect 792 991 862 1025
rect 896 991 902 1025
rect 792 953 902 991
rect 792 919 862 953
rect 896 919 902 953
rect 792 881 902 919
rect 792 847 862 881
rect 896 847 902 881
rect 792 809 902 847
rect 792 775 862 809
rect 896 775 902 809
rect 792 737 902 775
rect 792 703 862 737
rect 896 703 902 737
rect 792 665 902 703
rect 792 631 862 665
rect 896 631 902 665
rect 792 593 902 631
rect 792 559 862 593
rect 896 559 902 593
rect 792 521 902 559
rect 792 487 862 521
rect 896 487 902 521
rect 792 449 902 487
rect 792 415 862 449
rect 896 415 902 449
rect 792 377 902 415
rect 792 343 862 377
rect 896 343 902 377
rect 792 305 902 343
rect 792 271 862 305
rect 896 271 902 305
rect 792 233 902 271
rect 792 199 862 233
rect 896 199 902 233
rect 792 161 902 199
rect 792 127 862 161
rect 896 127 902 161
rect 792 89 902 127
rect 792 55 862 89
rect 896 55 902 89
rect 792 17 902 55
rect 792 -17 862 17
rect 896 -17 902 17
rect 792 -55 902 -17
rect 792 -89 862 -55
rect 896 -89 902 -55
rect 792 -127 902 -89
rect 792 -161 862 -127
rect 896 -161 902 -127
rect 792 -199 902 -161
rect 792 -233 862 -199
rect 896 -233 902 -199
rect 792 -271 902 -233
rect 792 -305 862 -271
rect 896 -305 902 -271
rect 792 -343 902 -305
rect 792 -377 862 -343
rect 896 -377 902 -343
rect 792 -415 902 -377
rect 792 -449 862 -415
rect 896 -449 902 -415
rect 792 -487 902 -449
rect 792 -521 862 -487
rect 896 -521 902 -487
rect 792 -559 902 -521
rect 792 -593 862 -559
rect 896 -593 902 -559
rect 792 -631 902 -593
rect 792 -665 862 -631
rect 896 -665 902 -631
rect 792 -703 902 -665
rect 792 -737 862 -703
rect 896 -737 902 -703
rect 792 -775 902 -737
rect 792 -809 862 -775
rect 896 -809 902 -775
rect 792 -847 902 -809
rect 792 -881 862 -847
rect 896 -881 902 -847
rect 792 -919 902 -881
rect 792 -953 862 -919
rect 896 -953 902 -919
rect 792 -991 902 -953
rect 792 -1025 862 -991
rect 896 -1025 902 -991
rect 792 -1063 902 -1025
rect 792 -1097 862 -1063
rect 896 -1097 902 -1063
rect 792 -1135 902 -1097
rect 792 -1169 862 -1135
rect 896 -1169 902 -1135
rect 792 -1207 902 -1169
rect 792 -1241 862 -1207
rect 896 -1241 902 -1207
rect 792 -1279 902 -1241
rect 792 -1313 862 -1279
rect 896 -1313 902 -1279
rect 792 -1351 902 -1313
rect 792 -1385 862 -1351
rect 896 -1385 902 -1351
rect 792 -1423 902 -1385
rect 792 -1457 862 -1423
rect 896 -1457 902 -1423
rect 792 -1495 902 -1457
rect 792 -1529 862 -1495
rect 896 -1529 902 -1495
rect 792 -1567 902 -1529
rect 792 -1601 862 -1567
rect 896 -1601 902 -1567
rect 792 -1639 902 -1601
rect 792 -1673 862 -1639
rect 896 -1673 902 -1639
rect 792 -1711 902 -1673
rect 792 -1745 862 -1711
rect 896 -1745 902 -1711
rect 792 -1783 902 -1745
rect 792 -1817 862 -1783
rect 896 -1817 902 -1783
rect 792 -1855 902 -1817
rect 792 -1889 862 -1855
rect 896 -1889 902 -1855
rect 792 -1927 902 -1889
rect 792 -1961 862 -1927
rect 896 -1961 902 -1927
rect 792 -1999 902 -1961
rect 792 -2033 862 -1999
rect 896 -2033 902 -1999
rect 792 -2071 902 -2033
rect 792 -2105 862 -2071
rect 896 -2105 902 -2071
rect 792 -2143 902 -2105
rect 792 -2177 862 -2143
rect 896 -2177 902 -2143
rect 792 -2215 902 -2177
rect 792 -2249 862 -2215
rect 896 -2249 902 -2215
rect 792 -2287 902 -2249
rect 792 -2321 862 -2287
rect 896 -2321 902 -2287
rect 792 -2359 902 -2321
rect 792 -2393 862 -2359
rect 896 -2393 902 -2359
rect 792 -2431 902 -2393
rect 792 -2465 862 -2431
rect 896 -2465 902 -2431
rect 792 -2503 902 -2465
rect 792 -2537 862 -2503
rect 896 -2537 902 -2503
rect 792 -2575 902 -2537
rect 792 -2609 862 -2575
rect 896 -2609 902 -2575
rect 792 -2647 902 -2609
rect 792 -2681 862 -2647
rect 896 -2681 902 -2647
rect 792 -2719 902 -2681
rect 792 -2753 862 -2719
rect 896 -2753 902 -2719
rect 792 -2791 902 -2753
rect 792 -2825 862 -2791
rect 896 -2825 902 -2791
rect 792 -2863 902 -2825
rect 792 -2897 862 -2863
rect 896 -2897 902 -2863
rect 792 -2935 902 -2897
rect 792 -2969 862 -2935
rect 896 -2969 902 -2935
rect 792 -3007 902 -2969
rect 792 -3041 862 -3007
rect 896 -3041 902 -3007
rect 792 -3079 902 -3041
rect 792 -3113 862 -3079
rect 896 -3113 902 -3079
rect 792 -3151 902 -3113
rect 792 -3185 862 -3151
rect 896 -3185 902 -3151
rect 792 -3223 902 -3185
rect 792 -3257 862 -3223
rect 896 -3257 902 -3223
rect 792 -3295 902 -3257
rect 792 -3329 862 -3295
rect 896 -3329 902 -3295
rect 792 -3367 902 -3329
rect 792 -3401 862 -3367
rect 896 -3401 902 -3367
rect 792 -3439 902 -3401
rect 792 -3473 862 -3439
rect 896 -3473 902 -3439
rect 792 -3511 902 -3473
rect 792 -3545 862 -3511
rect 896 -3545 902 -3511
rect 792 -3583 902 -3545
rect 792 -3617 862 -3583
rect 896 -3617 902 -3583
rect 792 -3655 902 -3617
rect 792 -3689 862 -3655
rect 896 -3689 902 -3655
rect 792 -3727 902 -3689
rect 792 -3761 862 -3727
rect 896 -3761 902 -3727
rect 792 -3799 902 -3761
rect 792 -3833 862 -3799
rect 896 -3833 902 -3799
rect 792 -3871 902 -3833
rect 792 -3905 862 -3871
rect 896 -3905 902 -3871
rect 792 -3943 902 -3905
rect 792 -3977 862 -3943
rect 896 -3977 902 -3943
rect 792 -4015 902 -3977
rect 792 -4049 862 -4015
rect 896 -4049 902 -4015
rect 792 -4087 902 -4049
rect 792 -4121 862 -4087
rect 896 -4121 902 -4087
rect 792 -4159 902 -4121
rect 792 -4193 862 -4159
rect 896 -4193 902 -4159
rect 792 -4231 902 -4193
rect 792 -4265 862 -4231
rect 896 -4265 902 -4231
rect 792 -4303 902 -4265
rect 792 -4337 862 -4303
rect 896 -4337 902 -4303
rect 792 -4375 902 -4337
rect 792 -4409 862 -4375
rect 896 -4409 902 -4375
rect 792 -4447 902 -4409
rect 792 -4481 862 -4447
rect 896 -4481 902 -4447
rect 792 -4519 902 -4481
rect 792 -4553 862 -4519
rect 896 -4553 902 -4519
rect 792 -4591 902 -4553
rect 792 -4625 862 -4591
rect 896 -4625 902 -4591
rect 792 -4663 902 -4625
rect 792 -4697 862 -4663
rect 896 -4697 902 -4663
rect 792 -4735 902 -4697
rect 792 -4769 862 -4735
rect 896 -4769 902 -4735
rect 792 -4807 902 -4769
rect 792 -4841 862 -4807
rect 896 -4841 902 -4807
rect 792 -4879 902 -4841
rect 792 -4913 862 -4879
rect 896 -4913 902 -4879
rect 792 -4951 902 -4913
rect 792 -4985 862 -4951
rect 896 -4985 902 -4951
rect 792 -5062 902 -4985
tri 970 5000 990 5020 se
rect 990 5000 1138 5020
tri 1138 5000 1158 5020 sw
rect 970 4985 1158 5000
rect 970 -4985 1011 4985
rect 1117 -4985 1158 4985
rect 970 -5000 1158 -4985
tri 970 -5020 990 -5000 ne
rect 990 -5020 1138 -5000
tri 1138 -5020 1158 -5000 nw
rect 1226 4985 1330 5062
rect 1226 4951 1232 4985
rect 1266 4951 1330 4985
rect 1226 4913 1330 4951
rect 1226 4879 1232 4913
rect 1266 4879 1330 4913
rect 1226 4841 1330 4879
rect 1226 4807 1232 4841
rect 1266 4807 1330 4841
rect 1226 4769 1330 4807
rect 1226 4735 1232 4769
rect 1266 4735 1330 4769
rect 1226 4697 1330 4735
rect 1226 4663 1232 4697
rect 1266 4663 1330 4697
rect 1226 4625 1330 4663
rect 1226 4591 1232 4625
rect 1266 4591 1330 4625
rect 1226 4553 1330 4591
rect 1226 4519 1232 4553
rect 1266 4519 1330 4553
rect 1226 4481 1330 4519
rect 1226 4447 1232 4481
rect 1266 4447 1330 4481
rect 1226 4409 1330 4447
rect 1226 4375 1232 4409
rect 1266 4375 1330 4409
rect 1226 4337 1330 4375
rect 1226 4303 1232 4337
rect 1266 4303 1330 4337
rect 1226 4265 1330 4303
rect 1226 4231 1232 4265
rect 1266 4231 1330 4265
rect 1226 4193 1330 4231
rect 1226 4159 1232 4193
rect 1266 4159 1330 4193
rect 1226 4121 1330 4159
rect 1226 4087 1232 4121
rect 1266 4087 1330 4121
rect 1226 4049 1330 4087
rect 1226 4015 1232 4049
rect 1266 4015 1330 4049
rect 1226 3977 1330 4015
rect 1226 3943 1232 3977
rect 1266 3943 1330 3977
rect 1226 3905 1330 3943
rect 1226 3871 1232 3905
rect 1266 3871 1330 3905
rect 1226 3833 1330 3871
rect 1226 3799 1232 3833
rect 1266 3799 1330 3833
rect 1226 3761 1330 3799
rect 1226 3727 1232 3761
rect 1266 3727 1330 3761
rect 1226 3689 1330 3727
rect 1226 3655 1232 3689
rect 1266 3655 1330 3689
rect 1226 3617 1330 3655
rect 1226 3583 1232 3617
rect 1266 3583 1330 3617
rect 1226 3545 1330 3583
rect 1226 3511 1232 3545
rect 1266 3511 1330 3545
rect 1226 3473 1330 3511
rect 1226 3439 1232 3473
rect 1266 3439 1330 3473
rect 1226 3401 1330 3439
rect 1226 3367 1232 3401
rect 1266 3367 1330 3401
rect 1226 3329 1330 3367
rect 1226 3295 1232 3329
rect 1266 3295 1330 3329
rect 1226 3257 1330 3295
rect 1226 3223 1232 3257
rect 1266 3223 1330 3257
rect 1226 3185 1330 3223
rect 1226 3151 1232 3185
rect 1266 3151 1330 3185
rect 1226 3113 1330 3151
rect 1226 3079 1232 3113
rect 1266 3079 1330 3113
rect 1226 3041 1330 3079
rect 1226 3007 1232 3041
rect 1266 3007 1330 3041
rect 1226 2969 1330 3007
rect 1226 2935 1232 2969
rect 1266 2935 1330 2969
rect 1226 2897 1330 2935
rect 1226 2863 1232 2897
rect 1266 2863 1330 2897
rect 1226 2825 1330 2863
rect 1226 2791 1232 2825
rect 1266 2791 1330 2825
rect 1226 2753 1330 2791
rect 1226 2719 1232 2753
rect 1266 2719 1330 2753
rect 1226 2681 1330 2719
rect 1226 2647 1232 2681
rect 1266 2647 1330 2681
rect 1226 2609 1330 2647
rect 1226 2575 1232 2609
rect 1266 2575 1330 2609
rect 1226 2537 1330 2575
rect 1226 2503 1232 2537
rect 1266 2503 1330 2537
rect 1226 2465 1330 2503
rect 1226 2431 1232 2465
rect 1266 2431 1330 2465
rect 1226 2393 1330 2431
rect 1226 2359 1232 2393
rect 1266 2359 1330 2393
rect 1226 2321 1330 2359
rect 1226 2287 1232 2321
rect 1266 2287 1330 2321
rect 1226 2249 1330 2287
rect 1226 2215 1232 2249
rect 1266 2215 1330 2249
rect 1226 2177 1330 2215
rect 1226 2143 1232 2177
rect 1266 2143 1330 2177
rect 1226 2105 1330 2143
rect 1226 2071 1232 2105
rect 1266 2071 1330 2105
rect 1226 2033 1330 2071
rect 1226 1999 1232 2033
rect 1266 1999 1330 2033
rect 1226 1961 1330 1999
rect 1226 1927 1232 1961
rect 1266 1927 1330 1961
rect 1226 1889 1330 1927
rect 1226 1855 1232 1889
rect 1266 1855 1330 1889
rect 1226 1817 1330 1855
rect 1226 1783 1232 1817
rect 1266 1783 1330 1817
rect 1226 1745 1330 1783
rect 1226 1711 1232 1745
rect 1266 1711 1330 1745
rect 1226 1673 1330 1711
rect 1226 1639 1232 1673
rect 1266 1639 1330 1673
rect 1226 1601 1330 1639
rect 1226 1567 1232 1601
rect 1266 1567 1330 1601
rect 1226 1529 1330 1567
rect 1226 1495 1232 1529
rect 1266 1495 1330 1529
rect 1226 1457 1330 1495
rect 1226 1423 1232 1457
rect 1266 1423 1330 1457
rect 1226 1385 1330 1423
rect 1226 1351 1232 1385
rect 1266 1351 1330 1385
rect 1226 1313 1330 1351
rect 1226 1279 1232 1313
rect 1266 1279 1330 1313
rect 1226 1241 1330 1279
rect 1226 1207 1232 1241
rect 1266 1207 1330 1241
rect 1226 1169 1330 1207
rect 1226 1135 1232 1169
rect 1266 1135 1330 1169
rect 1226 1097 1330 1135
rect 1226 1063 1232 1097
rect 1266 1063 1330 1097
rect 1226 1025 1330 1063
rect 1226 991 1232 1025
rect 1266 991 1330 1025
rect 1226 953 1330 991
rect 1226 919 1232 953
rect 1266 919 1330 953
rect 1226 881 1330 919
rect 1226 847 1232 881
rect 1266 847 1330 881
rect 1226 809 1330 847
rect 1226 775 1232 809
rect 1266 775 1330 809
rect 1226 737 1330 775
rect 1226 703 1232 737
rect 1266 703 1330 737
rect 1226 665 1330 703
rect 1226 631 1232 665
rect 1266 631 1330 665
rect 1226 593 1330 631
rect 1226 559 1232 593
rect 1266 559 1330 593
rect 1226 521 1330 559
rect 1226 487 1232 521
rect 1266 487 1330 521
rect 1226 449 1330 487
rect 1226 415 1232 449
rect 1266 415 1330 449
rect 1226 377 1330 415
rect 1226 343 1232 377
rect 1266 343 1330 377
rect 1226 305 1330 343
rect 1226 271 1232 305
rect 1266 271 1330 305
rect 1226 233 1330 271
rect 1226 199 1232 233
rect 1266 199 1330 233
rect 1226 161 1330 199
rect 1226 127 1232 161
rect 1266 127 1330 161
rect 1226 89 1330 127
rect 1226 55 1232 89
rect 1266 55 1330 89
rect 1226 17 1330 55
rect 1226 -17 1232 17
rect 1266 -17 1330 17
rect 1226 -55 1330 -17
rect 1226 -89 1232 -55
rect 1266 -89 1330 -55
rect 1226 -127 1330 -89
rect 1226 -161 1232 -127
rect 1266 -161 1330 -127
rect 1226 -199 1330 -161
rect 1226 -233 1232 -199
rect 1266 -233 1330 -199
rect 1226 -271 1330 -233
rect 1226 -305 1232 -271
rect 1266 -305 1330 -271
rect 1226 -343 1330 -305
rect 1226 -377 1232 -343
rect 1266 -377 1330 -343
rect 1226 -415 1330 -377
rect 1226 -449 1232 -415
rect 1266 -449 1330 -415
rect 1226 -487 1330 -449
rect 1226 -521 1232 -487
rect 1266 -521 1330 -487
rect 1226 -559 1330 -521
rect 1226 -593 1232 -559
rect 1266 -593 1330 -559
rect 1226 -631 1330 -593
rect 1226 -665 1232 -631
rect 1266 -665 1330 -631
rect 1226 -703 1330 -665
rect 1226 -737 1232 -703
rect 1266 -737 1330 -703
rect 1226 -775 1330 -737
rect 1226 -809 1232 -775
rect 1266 -809 1330 -775
rect 1226 -847 1330 -809
rect 1226 -881 1232 -847
rect 1266 -881 1330 -847
rect 1226 -919 1330 -881
rect 1226 -953 1232 -919
rect 1266 -953 1330 -919
rect 1226 -991 1330 -953
rect 1226 -1025 1232 -991
rect 1266 -1025 1330 -991
rect 1226 -1063 1330 -1025
rect 1226 -1097 1232 -1063
rect 1266 -1097 1330 -1063
rect 1226 -1135 1330 -1097
rect 1226 -1169 1232 -1135
rect 1266 -1169 1330 -1135
rect 1226 -1207 1330 -1169
rect 1226 -1241 1232 -1207
rect 1266 -1241 1330 -1207
rect 1226 -1279 1330 -1241
rect 1226 -1313 1232 -1279
rect 1266 -1313 1330 -1279
rect 1226 -1351 1330 -1313
rect 1226 -1385 1232 -1351
rect 1266 -1385 1330 -1351
rect 1226 -1423 1330 -1385
rect 1226 -1457 1232 -1423
rect 1266 -1457 1330 -1423
rect 1226 -1495 1330 -1457
rect 1226 -1529 1232 -1495
rect 1266 -1529 1330 -1495
rect 1226 -1567 1330 -1529
rect 1226 -1601 1232 -1567
rect 1266 -1601 1330 -1567
rect 1226 -1639 1330 -1601
rect 1226 -1673 1232 -1639
rect 1266 -1673 1330 -1639
rect 1226 -1711 1330 -1673
rect 1226 -1745 1232 -1711
rect 1266 -1745 1330 -1711
rect 1226 -1783 1330 -1745
rect 1226 -1817 1232 -1783
rect 1266 -1817 1330 -1783
rect 1226 -1855 1330 -1817
rect 1226 -1889 1232 -1855
rect 1266 -1889 1330 -1855
rect 1226 -1927 1330 -1889
rect 1226 -1961 1232 -1927
rect 1266 -1961 1330 -1927
rect 1226 -1999 1330 -1961
rect 1226 -2033 1232 -1999
rect 1266 -2033 1330 -1999
rect 1226 -2071 1330 -2033
rect 1226 -2105 1232 -2071
rect 1266 -2105 1330 -2071
rect 1226 -2143 1330 -2105
rect 1226 -2177 1232 -2143
rect 1266 -2177 1330 -2143
rect 1226 -2215 1330 -2177
rect 1226 -2249 1232 -2215
rect 1266 -2249 1330 -2215
rect 1226 -2287 1330 -2249
rect 1226 -2321 1232 -2287
rect 1266 -2321 1330 -2287
rect 1226 -2359 1330 -2321
rect 1226 -2393 1232 -2359
rect 1266 -2393 1330 -2359
rect 1226 -2431 1330 -2393
rect 1226 -2465 1232 -2431
rect 1266 -2465 1330 -2431
rect 1226 -2503 1330 -2465
rect 1226 -2537 1232 -2503
rect 1266 -2537 1330 -2503
rect 1226 -2575 1330 -2537
rect 1226 -2609 1232 -2575
rect 1266 -2609 1330 -2575
rect 1226 -2647 1330 -2609
rect 1226 -2681 1232 -2647
rect 1266 -2681 1330 -2647
rect 1226 -2719 1330 -2681
rect 1226 -2753 1232 -2719
rect 1266 -2753 1330 -2719
rect 1226 -2791 1330 -2753
rect 1226 -2825 1232 -2791
rect 1266 -2825 1330 -2791
rect 1226 -2863 1330 -2825
rect 1226 -2897 1232 -2863
rect 1266 -2897 1330 -2863
rect 1226 -2935 1330 -2897
rect 1226 -2969 1232 -2935
rect 1266 -2969 1330 -2935
rect 1226 -3007 1330 -2969
rect 1226 -3041 1232 -3007
rect 1266 -3041 1330 -3007
rect 1226 -3079 1330 -3041
rect 1226 -3113 1232 -3079
rect 1266 -3113 1330 -3079
rect 1226 -3151 1330 -3113
rect 1226 -3185 1232 -3151
rect 1266 -3185 1330 -3151
rect 1226 -3223 1330 -3185
rect 1226 -3257 1232 -3223
rect 1266 -3257 1330 -3223
rect 1226 -3295 1330 -3257
rect 1226 -3329 1232 -3295
rect 1266 -3329 1330 -3295
rect 1226 -3367 1330 -3329
rect 1226 -3401 1232 -3367
rect 1266 -3401 1330 -3367
rect 1226 -3439 1330 -3401
rect 1226 -3473 1232 -3439
rect 1266 -3473 1330 -3439
rect 1226 -3511 1330 -3473
rect 1226 -3545 1232 -3511
rect 1266 -3545 1330 -3511
rect 1226 -3583 1330 -3545
rect 1226 -3617 1232 -3583
rect 1266 -3617 1330 -3583
rect 1226 -3655 1330 -3617
rect 1226 -3689 1232 -3655
rect 1266 -3689 1330 -3655
rect 1226 -3727 1330 -3689
rect 1226 -3761 1232 -3727
rect 1266 -3761 1330 -3727
rect 1226 -3799 1330 -3761
rect 1226 -3833 1232 -3799
rect 1266 -3833 1330 -3799
rect 1226 -3871 1330 -3833
rect 1226 -3905 1232 -3871
rect 1266 -3905 1330 -3871
rect 1226 -3943 1330 -3905
rect 1226 -3977 1232 -3943
rect 1266 -3977 1330 -3943
rect 1226 -4015 1330 -3977
rect 1226 -4049 1232 -4015
rect 1266 -4049 1330 -4015
rect 1226 -4087 1330 -4049
rect 1226 -4121 1232 -4087
rect 1266 -4121 1330 -4087
rect 1226 -4159 1330 -4121
rect 1226 -4193 1232 -4159
rect 1266 -4193 1330 -4159
rect 1226 -4231 1330 -4193
rect 1226 -4265 1232 -4231
rect 1266 -4265 1330 -4231
rect 1226 -4303 1330 -4265
rect 1226 -4337 1232 -4303
rect 1266 -4337 1330 -4303
rect 1226 -4375 1330 -4337
rect 1226 -4409 1232 -4375
rect 1266 -4409 1330 -4375
rect 1226 -4447 1330 -4409
rect 1226 -4481 1232 -4447
rect 1266 -4481 1330 -4447
rect 1226 -4519 1330 -4481
rect 1226 -4553 1232 -4519
rect 1266 -4553 1330 -4519
rect 1226 -4591 1330 -4553
rect 1226 -4625 1232 -4591
rect 1266 -4625 1330 -4591
rect 1226 -4663 1330 -4625
rect 1226 -4697 1232 -4663
rect 1266 -4697 1330 -4663
rect 1226 -4735 1330 -4697
rect 1226 -4769 1232 -4735
rect 1266 -4769 1330 -4735
rect 1226 -4807 1330 -4769
rect 1226 -4841 1232 -4807
rect 1266 -4841 1330 -4807
rect 1226 -4879 1330 -4841
rect 1226 -4913 1232 -4879
rect 1266 -4913 1330 -4879
rect 1226 -4951 1330 -4913
rect 1226 -4985 1232 -4951
rect 1266 -4985 1330 -4951
tri 902 -5062 942 -5022 sw
tri 1186 -5062 1226 -5022 se
rect 1226 -5062 1330 -4985
rect 792 -5068 1330 -5062
rect 792 -5102 975 -5068
rect 1009 -5102 1047 -5068
rect 1081 -5102 1119 -5068
rect 1153 -5102 1330 -5068
rect 792 -5168 1330 -5102
rect 166 -5268 629 -5237
rect 1488 -5237 1542 5237
rect 1936 -5237 1956 5237
tri 629 -5268 651 -5246 sw
tri 1466 -5268 1488 -5246 se
rect 1488 -5268 1956 -5237
rect 166 -5286 651 -5268
tri 651 -5286 669 -5268 sw
tri 1448 -5286 1466 -5268 se
rect 1466 -5286 1956 -5268
rect 166 -5346 1956 -5286
rect 166 -5360 684 -5346
tri 166 -5740 546 -5360 ne
rect 546 -5740 684 -5360
rect 1438 -5360 1956 -5346
rect 1438 -5740 1556 -5360
tri 546 -5760 566 -5740 ne
rect 566 -5760 1556 -5740
tri 1556 -5760 1956 -5360 nw
<< properties >>
string FIXED_BBOX 879 -5085 1249 5085
string GDS_END 5160004
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io__analog.gds
string GDS_START 4824240
<< end >>
