magic
tech sky130A
magscale 1 2
timestamp 1681267127
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 1 21 624 203
rect 30 -17 64 21
<< locali >>
rect 288 401 354 493
rect 456 401 522 493
rect 288 367 522 401
rect 456 333 522 367
rect 456 299 627 333
rect 18 153 69 265
rect 173 199 248 265
rect 558 181 627 299
rect 288 147 627 181
rect 288 53 354 147
rect 456 53 522 147
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 31 333 103 493
rect 212 367 246 527
rect 388 435 422 527
rect 556 367 590 527
rect 31 299 323 333
rect 103 165 139 299
rect 282 249 323 299
rect 282 215 524 249
rect 21 17 69 119
rect 103 58 169 165
rect 212 17 246 165
rect 388 17 422 113
rect 556 17 590 113
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
rlabel locali s 173 199 248 265 6 A
port 1 nsew signal input
rlabel locali s 18 153 69 265 6 B
port 2 nsew signal input
rlabel metal1 s 0 -48 644 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 1 21 624 203 6 VNB
port 4 nsew ground bidirectional
rlabel nwell s -38 261 682 582 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 496 644 592 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 456 53 522 147 6 X
port 7 nsew signal output
rlabel locali s 288 53 354 147 6 X
port 7 nsew signal output
rlabel locali s 288 147 627 181 6 X
port 7 nsew signal output
rlabel locali s 558 181 627 299 6 X
port 7 nsew signal output
rlabel locali s 456 299 627 333 6 X
port 7 nsew signal output
rlabel locali s 456 333 522 367 6 X
port 7 nsew signal output
rlabel locali s 288 367 522 401 6 X
port 7 nsew signal output
rlabel locali s 456 401 522 493 6 X
port 7 nsew signal output
rlabel locali s 288 401 354 493 6 X
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 644 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 994424
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 988722
<< end >>
