magic
tech sky130A
magscale 1 2
timestamp 1681267127
use sky130_fd_pr__dfl1sd2__example_5595914180884  sky130_fd_pr__dfl1sd2__example_5595914180884_0
timestamp 1681267127
transform 1 0 120 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_5595914180884  sky130_fd_pr__dfl1sd2__example_5595914180884_1
timestamp 1681267127
transform 1 0 296 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_5595914180884  sky130_fd_pr__dfl1sd2__example_5595914180884_2
timestamp 1681267127
transform 1 0 472 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_5595914180884  sky130_fd_pr__dfl1sd2__example_5595914180884_3
timestamp 1681267127
transform 1 0 648 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_5595914180819  sky130_fd_pr__dfl1sd__example_5595914180819_0
timestamp 1681267127
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_5595914180819  sky130_fd_pr__dfl1sd__example_5595914180819_1
timestamp 1681267127
transform 1 0 824 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 7410124
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 7407146
<< end >>
