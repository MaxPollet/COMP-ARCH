magic
tech sky130A
magscale 1 2
timestamp 1681267127
<< nwell >>
rect -38 261 2706 582
<< pwell >>
rect 1408 157 1759 201
rect 2198 157 2667 203
rect 1 21 2667 157
rect 30 -17 64 21
<< locali >>
rect 17 153 69 335
rect 211 153 267 335
rect 581 318 617 392
rect 581 211 713 318
rect 581 145 620 211
rect 2300 51 2366 493
rect 2583 299 2651 490
rect 2614 165 2651 299
rect 2583 55 2651 165
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2668 561
rect 17 405 69 493
rect 103 439 153 527
rect 187 451 409 493
rect 187 405 221 451
rect 454 417 504 493
rect 538 428 606 527
rect 17 369 221 405
rect 259 374 339 415
rect 109 255 165 335
rect 109 221 122 255
rect 156 221 165 255
rect 109 153 165 221
rect 301 141 339 374
rect 373 354 504 417
rect 373 181 440 354
rect 474 255 540 320
rect 474 221 489 255
rect 523 221 540 255
rect 474 215 540 221
rect 651 391 685 465
rect 719 455 785 527
rect 819 427 888 493
rect 651 355 799 391
rect 373 143 503 181
rect 747 177 799 355
rect 299 133 339 141
rect 295 131 339 133
rect 295 129 334 131
rect 292 127 334 129
rect 289 126 334 127
rect 288 124 334 126
rect 286 123 334 124
rect 284 122 332 123
rect 281 121 332 122
rect 279 120 332 121
rect 17 17 96 119
rect 276 118 332 120
rect 276 112 331 118
rect 175 56 331 112
rect 365 17 401 109
rect 452 51 503 143
rect 654 143 799 177
rect 833 284 888 427
rect 922 323 966 493
rect 1006 427 1151 493
rect 1189 455 1255 527
rect 922 318 983 323
rect 932 289 983 318
rect 1041 315 1083 391
rect 833 218 898 284
rect 538 17 606 111
rect 654 51 691 143
rect 833 117 867 218
rect 932 184 966 289
rect 1117 279 1151 427
rect 1310 421 1353 490
rect 1401 425 1592 527
rect 1626 425 1787 492
rect 1839 447 1905 527
rect 1185 387 1353 421
rect 1753 413 1787 425
rect 1939 413 1982 490
rect 2027 447 2093 527
rect 1185 315 1219 387
rect 1328 289 1403 353
rect 1438 299 1601 391
rect 1017 255 1287 279
rect 1460 255 1532 265
rect 726 17 788 109
rect 822 51 867 117
rect 901 51 966 184
rect 1000 245 1532 255
rect 1000 51 1088 245
rect 1122 161 1195 203
rect 1250 195 1532 245
rect 1567 179 1601 299
rect 1673 215 1719 381
rect 1753 379 2093 413
rect 1777 323 2015 345
rect 1811 305 2015 323
rect 2049 305 2093 379
rect 1811 289 1822 305
rect 1777 283 1822 289
rect 2127 271 2179 493
rect 2224 297 2266 527
rect 1762 179 1808 249
rect 1122 127 1307 161
rect 1122 17 1219 93
rect 1255 51 1307 127
rect 1347 17 1526 161
rect 1567 139 1808 179
rect 1858 237 2179 271
rect 1858 171 1893 237
rect 1931 169 2109 203
rect 1931 89 1965 169
rect 1682 55 1965 89
rect 2044 17 2078 109
rect 2143 108 2179 237
rect 2112 51 2179 108
rect 2224 17 2266 177
rect 2412 265 2454 493
rect 2515 315 2549 527
rect 2412 199 2580 265
rect 2412 51 2454 199
rect 2508 17 2549 165
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2668 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 2513 527 2547 561
rect 2605 527 2639 561
rect 122 221 156 255
rect 489 221 523 255
rect 1777 289 1811 323
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
rect 2513 -17 2547 17
rect 2605 -17 2639 17
<< metal1 >>
rect 0 561 2668 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2668 561
rect 0 496 2668 527
rect 1316 320 1374 329
rect 1765 323 1823 329
rect 1765 320 1777 323
rect 1316 292 1777 320
rect 1316 283 1374 292
rect 1765 289 1777 292
rect 1811 289 1823 323
rect 1765 283 1823 289
rect 110 255 168 261
rect 110 221 122 255
rect 156 252 168 255
rect 477 255 535 261
rect 477 252 489 255
rect 156 224 489 252
rect 156 221 168 224
rect 110 215 168 221
rect 477 221 489 224
rect 523 221 535 255
rect 477 215 535 221
rect 0 17 2668 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2668 17
rect 0 -48 2668 -17
<< obsm1 >>
rect 753 388 811 397
rect 1029 388 1087 397
rect 1489 388 1547 397
rect 753 360 1547 388
rect 753 351 811 360
rect 1029 351 1087 360
rect 1489 351 1547 360
rect 293 320 351 329
rect 937 320 995 329
rect 293 292 995 320
rect 293 283 351 292
rect 937 283 995 292
rect 845 252 903 261
rect 1673 252 1731 261
rect 845 224 1731 252
rect 845 215 903 224
rect 1673 215 1731 224
<< labels >>
rlabel locali s 581 145 620 211 6 CLK
port 1 nsew clock input
rlabel locali s 581 211 713 318 6 CLK
port 1 nsew clock input
rlabel locali s 581 318 617 392 6 CLK
port 1 nsew clock input
rlabel locali s 211 153 267 335 6 D
port 2 nsew signal input
rlabel locali s 17 153 69 335 6 SCD
port 3 nsew signal input
rlabel metal1 s 477 215 535 224 6 SCE
port 4 nsew signal input
rlabel metal1 s 110 215 168 224 6 SCE
port 4 nsew signal input
rlabel metal1 s 110 224 535 252 6 SCE
port 4 nsew signal input
rlabel metal1 s 477 252 535 261 6 SCE
port 4 nsew signal input
rlabel metal1 s 110 252 168 261 6 SCE
port 4 nsew signal input
rlabel metal1 s 1765 283 1823 292 6 SET_B
port 5 nsew signal input
rlabel metal1 s 1316 283 1374 292 6 SET_B
port 5 nsew signal input
rlabel metal1 s 1316 292 1823 320 6 SET_B
port 5 nsew signal input
rlabel metal1 s 1765 320 1823 329 6 SET_B
port 5 nsew signal input
rlabel metal1 s 1316 320 1374 329 6 SET_B
port 5 nsew signal input
rlabel metal1 s 0 -48 2668 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 1 21 2667 157 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 2198 157 2667 203 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 1408 157 1759 201 6 VNB
port 7 nsew ground bidirectional
rlabel nwell s -38 261 2706 582 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 496 2668 592 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 2583 55 2651 165 6 Q
port 10 nsew signal output
rlabel locali s 2614 165 2651 299 6 Q
port 10 nsew signal output
rlabel locali s 2583 299 2651 490 6 Q
port 10 nsew signal output
rlabel locali s 2300 51 2366 493 6 Q_N
port 11 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 2668 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 53504
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 31832
<< end >>
