magic
tech sky130A
magscale 1 2
timestamp 1681267127
<< nwell >>
rect -66 377 738 897
<< pwell >>
rect 50 43 668 283
rect -26 -43 698 43
<< mvnmos >>
rect 133 107 233 257
rect 289 107 389 257
rect 489 173 589 257
<< mvpmos >>
rect 129 443 229 743
rect 285 443 385 743
rect 485 443 585 593
<< mvndiff >>
rect 76 249 133 257
rect 76 215 88 249
rect 122 215 133 249
rect 76 149 133 215
rect 76 115 88 149
rect 122 115 133 149
rect 76 107 133 115
rect 233 249 289 257
rect 233 215 244 249
rect 278 215 289 249
rect 233 149 289 215
rect 233 115 244 149
rect 278 115 289 149
rect 233 107 289 115
rect 389 249 489 257
rect 389 215 400 249
rect 434 215 489 249
rect 389 173 489 215
rect 589 232 642 257
rect 589 198 600 232
rect 634 198 642 232
rect 589 173 642 198
rect 389 149 446 173
rect 389 115 400 149
rect 434 115 446 149
rect 389 107 446 115
<< mvpdiff >>
rect 72 735 129 743
rect 72 701 84 735
rect 118 701 129 735
rect 72 652 129 701
rect 72 618 84 652
rect 118 618 129 652
rect 72 568 129 618
rect 72 534 84 568
rect 118 534 129 568
rect 72 485 129 534
rect 72 451 84 485
rect 118 451 129 485
rect 72 443 129 451
rect 229 735 285 743
rect 229 701 240 735
rect 274 701 285 735
rect 229 652 285 701
rect 229 618 240 652
rect 274 618 285 652
rect 229 568 285 618
rect 229 534 240 568
rect 274 534 285 568
rect 229 485 285 534
rect 229 451 240 485
rect 274 451 285 485
rect 229 443 285 451
rect 385 735 442 743
rect 385 701 396 735
rect 430 701 442 735
rect 385 655 442 701
rect 385 621 396 655
rect 430 621 442 655
rect 385 593 442 621
rect 385 574 485 593
rect 385 540 396 574
rect 430 540 485 574
rect 385 494 485 540
rect 385 460 396 494
rect 430 460 485 494
rect 385 443 485 460
rect 585 585 642 593
rect 585 551 596 585
rect 630 551 642 585
rect 585 485 642 551
rect 585 451 596 485
rect 630 451 642 485
rect 585 443 642 451
<< mvndiffc >>
rect 88 215 122 249
rect 88 115 122 149
rect 244 215 278 249
rect 244 115 278 149
rect 400 215 434 249
rect 600 198 634 232
rect 400 115 434 149
<< mvpdiffc >>
rect 84 701 118 735
rect 84 618 118 652
rect 84 534 118 568
rect 84 451 118 485
rect 240 701 274 735
rect 240 618 274 652
rect 240 534 274 568
rect 240 451 274 485
rect 396 701 430 735
rect 396 621 430 655
rect 396 540 430 574
rect 396 460 430 494
rect 596 551 630 585
rect 596 451 630 485
<< mvpsubdiff >>
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< mvnsubdiff >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 672 831
<< mvpsubdiffcont >>
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< mvnsubdiffcont >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
<< poly >>
rect 129 421 229 443
rect 129 379 233 421
rect 285 379 385 443
rect 485 421 585 443
rect 485 395 589 421
rect 129 335 389 379
rect 129 301 326 335
rect 360 301 389 335
rect 129 279 389 301
rect 485 361 505 395
rect 539 361 589 395
rect 485 279 589 361
rect 133 257 233 279
rect 289 257 389 279
rect 489 257 589 279
<< polycont >>
rect 326 301 360 335
rect 505 361 539 395
<< locali >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 672 831
rect 18 735 204 751
rect 18 701 22 735
rect 56 701 84 735
rect 128 701 166 735
rect 200 701 204 735
rect 18 652 204 701
rect 18 618 84 652
rect 118 618 204 652
rect 18 568 204 618
rect 18 534 84 568
rect 118 534 204 568
rect 18 485 204 534
rect 18 451 84 485
rect 118 451 204 485
rect 18 435 204 451
rect 240 735 274 751
rect 240 652 274 701
rect 240 568 274 618
rect 240 485 274 534
rect 310 735 560 751
rect 344 701 382 735
rect 430 701 454 735
rect 488 701 526 735
rect 310 655 560 701
rect 310 621 396 655
rect 430 621 560 655
rect 310 574 560 621
rect 310 540 396 574
rect 430 540 560 574
rect 310 494 560 540
rect 310 460 396 494
rect 430 460 560 494
rect 596 585 650 601
rect 630 551 650 585
rect 596 485 650 551
rect 240 356 274 451
rect 630 451 650 485
rect 25 344 274 356
rect 409 395 555 424
rect 409 361 505 395
rect 539 361 555 395
rect 409 355 555 361
rect 25 310 278 344
rect 18 249 208 265
rect 18 215 88 249
rect 122 215 208 249
rect 18 149 208 215
rect 18 115 88 149
rect 122 115 208 149
rect 18 113 208 115
rect 18 79 24 113
rect 58 79 96 113
rect 130 79 168 113
rect 202 79 208 113
rect 244 249 278 310
rect 314 335 373 351
rect 314 301 326 335
rect 360 319 373 335
rect 596 319 650 451
rect 360 301 650 319
rect 314 285 650 301
rect 244 149 278 215
rect 244 99 278 115
rect 314 215 400 249
rect 434 215 564 249
rect 314 149 564 215
rect 600 232 650 285
rect 634 198 650 232
rect 600 165 650 198
rect 314 115 400 149
rect 434 115 564 149
rect 314 113 564 115
rect 18 73 208 79
rect 348 79 386 113
rect 420 79 458 113
rect 492 79 530 113
rect 314 73 564 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 22 701 56 735
rect 94 701 118 735
rect 118 701 128 735
rect 166 701 200 735
rect 310 701 344 735
rect 382 701 396 735
rect 396 701 416 735
rect 454 701 488 735
rect 526 701 560 735
rect 24 79 58 113
rect 96 79 130 113
rect 168 79 202 113
rect 314 79 348 113
rect 386 79 420 113
rect 458 79 492 113
rect 530 79 564 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 831 672 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 672 831
rect 0 791 672 797
rect 0 735 672 763
rect 0 701 22 735
rect 56 701 94 735
rect 128 701 166 735
rect 200 701 310 735
rect 344 701 382 735
rect 416 701 454 735
rect 488 701 526 735
rect 560 701 672 735
rect 0 689 672 701
rect 0 113 672 125
rect 0 79 24 113
rect 58 79 96 113
rect 130 79 168 113
rect 202 79 314 113
rect 348 79 386 113
rect 420 79 458 113
rect 492 79 530 113
rect 564 79 672 113
rect 0 51 672 79
rect 0 17 672 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -23 672 -17
<< labels >>
rlabel comment s 0 0 0 0 4 buf_2
flabel metal1 s 0 51 672 125 0 FreeSans 340 0 0 0 VGND
port 2 nsew ground bidirectional
flabel metal1 s 0 0 672 23 0 FreeSans 340 0 0 0 VNB
port 3 nsew ground bidirectional
flabel metal1 s 0 689 672 763 0 FreeSans 340 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal1 s 0 791 672 814 0 FreeSans 340 0 0 0 VPB
port 4 nsew power bidirectional
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 672 814
string GDS_END 829860
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 821298
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
<< end >>
