magic
tech sky130A
timestamp 1681267127
<< properties >>
string GDS_END 30710716
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 30710012
<< end >>
