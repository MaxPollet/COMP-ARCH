magic
tech sky130A
magscale 1 2
timestamp 1681267127
<< nwell >>
rect -38 261 590 582
<< pwell >>
rect 1 21 545 203
rect 29 -17 63 21
<< locali >>
rect 121 265 155 450
rect 189 409 255 489
rect 395 409 535 493
rect 189 363 535 409
rect 189 319 255 363
rect 294 265 359 323
rect 17 199 79 265
rect 121 199 196 265
rect 260 199 359 265
rect 394 215 460 323
rect 494 169 535 363
rect 393 51 535 169
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 19 315 85 527
rect 289 455 355 527
rect 19 123 291 165
rect 19 51 85 123
rect 119 17 185 89
rect 225 51 291 123
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
<< metal1 >>
rect 0 561 552 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 0 496 552 527
rect 0 17 552 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
rect 0 -48 552 -17
<< labels >>
rlabel locali s 17 199 79 265 6 A1
port 1 nsew signal input
rlabel locali s 121 199 196 265 6 A2
port 2 nsew signal input
rlabel locali s 121 265 155 450 6 A2
port 2 nsew signal input
rlabel locali s 260 199 359 265 6 B1
port 3 nsew signal input
rlabel locali s 294 265 359 323 6 B1
port 3 nsew signal input
rlabel locali s 394 215 460 323 6 C1
port 4 nsew signal input
rlabel metal1 s 0 -48 552 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1 21 545 203 6 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 590 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 552 592 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 393 51 535 169 6 Y
port 9 nsew signal output
rlabel locali s 494 169 535 363 6 Y
port 9 nsew signal output
rlabel locali s 189 319 255 363 6 Y
port 9 nsew signal output
rlabel locali s 189 363 535 409 6 Y
port 9 nsew signal output
rlabel locali s 395 409 535 493 6 Y
port 9 nsew signal output
rlabel locali s 189 409 255 489 6 Y
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 552 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 776350
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 770954
<< end >>
