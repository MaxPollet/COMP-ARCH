magic
tech sky130A
magscale 1 2
timestamp 1681267127
use sky130_fd_pr__dfm1sd__example_55959141808169  sky130_fd_pr__dfm1sd__example_55959141808169_0
timestamp 1681267127
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfm1sd__example_55959141808169  sky130_fd_pr__dfm1sd__example_55959141808169_1
timestamp 1681267127
transform 1 0 100 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 39456338
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 39455288
<< end >>
