magic
tech sky130A
magscale 1 2
timestamp 1681267127
use sky130_fd_pr__hvdfl1sd__example_55959141808122  sky130_fd_pr__hvdfl1sd__example_55959141808122_0
timestamp 1681267127
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808122  sky130_fd_pr__hvdfl1sd__example_55959141808122_1
timestamp 1681267127
transform 1 0 200 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 39959788
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 39958734
<< end >>
