magic
tech sky130A
magscale 1 2
timestamp 1681267127
use sky130_fd_pr__dfl1sd2__example_55959141808679  sky130_fd_pr__dfl1sd2__example_55959141808679_0
timestamp 1681267127
transform 1 0 100 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808679  sky130_fd_pr__dfl1sd2__example_55959141808679_1
timestamp 1681267127
transform 1 0 256 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808679  sky130_fd_pr__dfl1sd2__example_55959141808679_2
timestamp 1681267127
transform 1 0 412 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808679  sky130_fd_pr__dfl1sd2__example_55959141808679_3
timestamp 1681267127
transform 1 0 568 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808679  sky130_fd_pr__dfl1sd2__example_55959141808679_4
timestamp 1681267127
transform 1 0 724 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808679  sky130_fd_pr__dfl1sd2__example_55959141808679_5
timestamp 1681267127
transform 1 0 880 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808679  sky130_fd_pr__dfl1sd2__example_55959141808679_6
timestamp 1681267127
transform 1 0 1036 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808679  sky130_fd_pr__dfl1sd2__example_55959141808679_7
timestamp 1681267127
transform 1 0 1192 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808679  sky130_fd_pr__dfl1sd2__example_55959141808679_8
timestamp 1681267127
transform 1 0 1348 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808679  sky130_fd_pr__dfl1sd2__example_55959141808679_9
timestamp 1681267127
transform 1 0 1504 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808679  sky130_fd_pr__dfl1sd2__example_55959141808679_10
timestamp 1681267127
transform 1 0 1660 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808679  sky130_fd_pr__dfl1sd2__example_55959141808679_11
timestamp 1681267127
transform 1 0 1816 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808679  sky130_fd_pr__dfl1sd2__example_55959141808679_12
timestamp 1681267127
transform 1 0 1972 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808679  sky130_fd_pr__dfl1sd2__example_55959141808679_13
timestamp 1681267127
transform 1 0 2128 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_55959141808678  sky130_fd_pr__dfl1sd__example_55959141808678_0
timestamp 1681267127
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_55959141808678  sky130_fd_pr__dfl1sd__example_55959141808678_1
timestamp 1681267127
transform 1 0 2284 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 11328814
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 11320668
<< end >>
