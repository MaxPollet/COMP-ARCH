magic
tech sky130A
magscale 1 2
timestamp 1681267127
<< nwell >>
rect -38 261 1602 582
<< pwell >>
rect 18 21 1561 203
rect 29 -17 63 21
<< scnmos >>
rect 97 47 127 177
rect 183 47 213 177
rect 269 47 299 177
rect 362 47 392 177
rect 459 47 489 177
rect 653 47 683 177
rect 740 47 770 177
rect 826 47 856 177
rect 1022 47 1052 177
rect 1108 47 1138 177
rect 1194 47 1224 177
rect 1280 47 1310 177
rect 1366 47 1396 177
rect 1452 47 1482 177
<< scpmoshvt >>
rect 83 297 113 497
rect 169 297 199 497
rect 255 297 285 497
rect 341 297 371 497
rect 529 297 559 497
rect 615 297 645 497
rect 748 297 778 497
rect 834 297 864 497
rect 1022 297 1052 497
rect 1108 297 1138 497
rect 1194 297 1224 497
rect 1280 297 1310 497
rect 1366 297 1396 497
rect 1452 297 1482 497
<< ndiff >>
rect 44 101 97 177
rect 44 67 52 101
rect 86 67 97 101
rect 44 47 97 67
rect 127 93 183 177
rect 127 59 138 93
rect 172 59 183 93
rect 127 47 183 59
rect 213 101 269 177
rect 213 67 224 101
rect 258 67 269 101
rect 213 47 269 67
rect 299 89 362 177
rect 299 55 318 89
rect 352 55 362 89
rect 299 47 362 55
rect 392 101 459 177
rect 392 67 403 101
rect 437 67 459 101
rect 392 47 459 67
rect 489 89 653 177
rect 489 55 500 89
rect 534 55 604 89
rect 638 55 653 89
rect 489 47 653 55
rect 683 169 740 177
rect 683 135 695 169
rect 729 135 740 169
rect 683 101 740 135
rect 683 67 695 101
rect 729 67 740 101
rect 683 47 740 67
rect 770 157 826 177
rect 770 123 781 157
rect 815 123 826 157
rect 770 47 826 123
rect 856 89 912 177
rect 856 55 866 89
rect 900 55 912 89
rect 856 47 912 55
rect 966 89 1022 177
rect 966 55 978 89
rect 1012 55 1022 89
rect 966 47 1022 55
rect 1052 101 1108 177
rect 1052 67 1063 101
rect 1097 67 1108 101
rect 1052 47 1108 67
rect 1138 89 1194 177
rect 1138 55 1149 89
rect 1183 55 1194 89
rect 1138 47 1194 55
rect 1224 101 1280 177
rect 1224 67 1235 101
rect 1269 67 1280 101
rect 1224 47 1280 67
rect 1310 89 1366 177
rect 1310 55 1321 89
rect 1355 55 1366 89
rect 1310 47 1366 55
rect 1396 101 1452 177
rect 1396 67 1407 101
rect 1441 67 1452 101
rect 1396 47 1452 67
rect 1482 93 1535 177
rect 1482 59 1493 93
rect 1527 59 1535 93
rect 1482 47 1535 59
<< pdiff >>
rect 30 477 83 497
rect 30 443 38 477
rect 72 443 83 477
rect 30 409 83 443
rect 30 375 38 409
rect 72 375 83 409
rect 30 297 83 375
rect 113 419 169 497
rect 113 385 124 419
rect 158 385 169 419
rect 113 351 169 385
rect 113 317 124 351
rect 158 317 169 351
rect 113 297 169 317
rect 199 477 255 497
rect 199 443 210 477
rect 244 443 255 477
rect 199 409 255 443
rect 199 375 210 409
rect 244 375 255 409
rect 199 341 255 375
rect 199 307 210 341
rect 244 307 255 341
rect 199 297 255 307
rect 285 419 341 497
rect 285 385 296 419
rect 330 385 341 419
rect 285 351 341 385
rect 285 317 296 351
rect 330 317 341 351
rect 285 297 341 317
rect 371 477 423 497
rect 371 443 381 477
rect 415 443 423 477
rect 371 409 423 443
rect 371 375 381 409
rect 415 375 423 409
rect 371 297 423 375
rect 477 467 529 497
rect 477 433 485 467
rect 519 433 529 467
rect 477 393 529 433
rect 477 359 485 393
rect 519 359 529 393
rect 477 297 529 359
rect 559 409 615 497
rect 559 375 570 409
rect 604 375 615 409
rect 559 341 615 375
rect 559 307 570 341
rect 604 307 615 341
rect 559 297 615 307
rect 645 465 748 497
rect 645 431 680 465
rect 714 431 748 465
rect 645 397 748 431
rect 645 363 680 397
rect 714 363 748 397
rect 645 297 748 363
rect 778 467 834 497
rect 778 433 789 467
rect 823 433 834 467
rect 778 297 834 433
rect 864 467 916 497
rect 864 433 874 467
rect 908 433 916 467
rect 864 399 916 433
rect 864 365 874 399
rect 908 365 916 399
rect 864 297 916 365
rect 970 485 1022 497
rect 970 451 978 485
rect 1012 451 1022 485
rect 970 297 1022 451
rect 1052 477 1108 497
rect 1052 443 1063 477
rect 1097 443 1108 477
rect 1052 409 1108 443
rect 1052 375 1063 409
rect 1097 375 1108 409
rect 1052 297 1108 375
rect 1138 485 1194 497
rect 1138 451 1149 485
rect 1183 451 1194 485
rect 1138 394 1194 451
rect 1138 360 1149 394
rect 1183 360 1194 394
rect 1138 297 1194 360
rect 1224 477 1280 497
rect 1224 443 1235 477
rect 1269 443 1280 477
rect 1224 384 1280 443
rect 1224 350 1235 384
rect 1269 350 1280 384
rect 1224 297 1280 350
rect 1310 485 1366 497
rect 1310 451 1321 485
rect 1355 451 1366 485
rect 1310 411 1366 451
rect 1310 377 1321 411
rect 1355 377 1366 411
rect 1310 297 1366 377
rect 1396 477 1452 497
rect 1396 443 1407 477
rect 1441 443 1452 477
rect 1396 384 1452 443
rect 1396 350 1407 384
rect 1441 350 1452 384
rect 1396 297 1452 350
rect 1482 485 1535 497
rect 1482 451 1493 485
rect 1527 451 1535 485
rect 1482 411 1535 451
rect 1482 377 1493 411
rect 1527 377 1535 411
rect 1482 297 1535 377
<< ndiffc >>
rect 52 67 86 101
rect 138 59 172 93
rect 224 67 258 101
rect 318 55 352 89
rect 403 67 437 101
rect 500 55 534 89
rect 604 55 638 89
rect 695 135 729 169
rect 695 67 729 101
rect 781 123 815 157
rect 866 55 900 89
rect 978 55 1012 89
rect 1063 67 1097 101
rect 1149 55 1183 89
rect 1235 67 1269 101
rect 1321 55 1355 89
rect 1407 67 1441 101
rect 1493 59 1527 93
<< pdiffc >>
rect 38 443 72 477
rect 38 375 72 409
rect 124 385 158 419
rect 124 317 158 351
rect 210 443 244 477
rect 210 375 244 409
rect 210 307 244 341
rect 296 385 330 419
rect 296 317 330 351
rect 381 443 415 477
rect 381 375 415 409
rect 485 433 519 467
rect 485 359 519 393
rect 570 375 604 409
rect 570 307 604 341
rect 680 431 714 465
rect 680 363 714 397
rect 789 433 823 467
rect 874 433 908 467
rect 874 365 908 399
rect 978 451 1012 485
rect 1063 443 1097 477
rect 1063 375 1097 409
rect 1149 451 1183 485
rect 1149 360 1183 394
rect 1235 443 1269 477
rect 1235 350 1269 384
rect 1321 451 1355 485
rect 1321 377 1355 411
rect 1407 443 1441 477
rect 1407 350 1441 384
rect 1493 451 1527 485
rect 1493 377 1527 411
<< poly >>
rect 21 249 199 265
rect 21 215 37 249
rect 71 215 199 249
rect 21 199 199 215
rect 255 249 403 264
rect 255 215 285 249
rect 319 215 353 249
rect 387 215 403 249
rect 255 199 403 215
rect 459 249 683 264
rect 459 215 506 249
rect 540 215 601 249
rect 635 215 683 249
rect 459 199 683 215
rect 740 249 899 267
rect 1022 259 1138 265
rect 740 215 781 249
rect 815 215 849 249
rect 883 215 899 249
rect 740 199 899 215
rect 991 249 1138 259
rect 991 215 1007 249
rect 1041 215 1075 249
rect 1109 215 1138 249
rect 991 205 1138 215
rect 1022 199 1138 205
rect 1194 249 1482 265
rect 1194 215 1210 249
rect 1244 215 1278 249
rect 1312 215 1346 249
rect 1380 215 1414 249
rect 1448 215 1482 249
rect 1194 199 1482 215
<< polycont >>
rect 37 215 71 249
rect 285 215 319 249
rect 353 215 387 249
rect 506 215 540 249
rect 601 215 635 249
rect 781 215 815 249
rect 849 215 883 249
rect 1007 215 1041 249
rect 1075 215 1109 249
rect 1210 215 1244 249
rect 1278 215 1312 249
rect 1346 215 1380 249
rect 1414 215 1448 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 22 477 432 493
rect 22 443 38 477
rect 72 459 210 477
rect 72 443 74 459
rect 22 409 74 443
rect 208 443 210 459
rect 244 459 381 477
rect 244 443 246 459
rect 22 375 38 409
rect 72 375 74 409
rect 22 359 74 375
rect 108 419 174 425
rect 108 385 124 419
rect 158 385 174 419
rect 108 351 174 385
rect 17 249 74 325
rect 17 215 37 249
rect 71 215 74 249
rect 17 195 74 215
rect 108 317 124 351
rect 158 317 174 351
rect 108 161 174 317
rect 208 409 246 443
rect 380 443 381 459
rect 415 443 432 477
rect 208 375 210 409
rect 244 375 246 409
rect 208 341 246 375
rect 208 307 210 341
rect 244 307 246 341
rect 208 291 246 307
rect 280 419 346 425
rect 280 385 296 419
rect 330 385 346 419
rect 280 351 346 385
rect 380 409 432 443
rect 380 375 381 409
rect 415 375 432 409
rect 380 359 432 375
rect 468 467 730 493
rect 468 433 485 467
rect 519 465 730 467
rect 519 459 680 465
rect 519 433 535 459
rect 468 393 535 433
rect 664 431 680 459
rect 714 431 730 465
rect 773 467 839 527
rect 961 485 1028 527
rect 773 433 789 467
rect 823 433 839 467
rect 873 467 925 483
rect 873 433 874 467
rect 908 433 925 467
rect 961 451 978 485
rect 1012 451 1028 485
rect 1062 477 1099 493
rect 468 359 485 393
rect 519 359 535 393
rect 569 409 620 425
rect 569 375 570 409
rect 604 375 620 409
rect 280 317 296 351
rect 330 325 346 351
rect 569 341 620 375
rect 664 399 730 431
rect 873 399 925 433
rect 1062 443 1063 477
rect 1097 443 1099 477
rect 1062 409 1099 443
rect 1062 399 1063 409
rect 664 397 874 399
rect 664 363 680 397
rect 714 365 874 397
rect 908 375 1063 399
rect 1097 375 1099 409
rect 908 365 1099 375
rect 714 363 1099 365
rect 664 359 1099 363
rect 1133 485 1199 527
rect 1133 451 1149 485
rect 1183 451 1199 485
rect 1133 394 1199 451
rect 1133 360 1149 394
rect 1183 360 1199 394
rect 1233 477 1271 493
rect 1233 443 1235 477
rect 1269 443 1271 477
rect 1233 384 1271 443
rect 569 325 570 341
rect 330 317 570 325
rect 280 307 570 317
rect 604 307 620 341
rect 1233 350 1235 384
rect 1269 350 1271 384
rect 1305 485 1371 527
rect 1305 451 1321 485
rect 1355 451 1371 485
rect 1305 411 1371 451
rect 1305 377 1321 411
rect 1355 377 1371 411
rect 1405 477 1443 493
rect 1405 443 1407 477
rect 1441 443 1443 477
rect 1405 384 1443 443
rect 1233 343 1271 350
rect 1405 350 1407 384
rect 1441 350 1443 384
rect 1477 485 1543 527
rect 1477 451 1493 485
rect 1527 451 1543 485
rect 1477 411 1543 451
rect 1477 377 1493 411
rect 1527 377 1543 411
rect 1477 361 1543 377
rect 1405 343 1443 350
rect 1233 327 1443 343
rect 280 291 620 307
rect 693 289 1195 325
rect 1233 293 1547 327
rect 208 249 456 257
rect 208 215 285 249
rect 319 215 353 249
rect 387 215 456 249
rect 208 195 456 215
rect 490 249 651 257
rect 490 215 506 249
rect 540 215 601 249
rect 635 215 651 249
rect 490 195 651 215
rect 693 169 731 289
rect 765 249 899 255
rect 765 215 781 249
rect 815 215 849 249
rect 883 215 899 249
rect 935 249 1125 255
rect 935 215 1007 249
rect 1041 215 1075 249
rect 1109 215 1125 249
rect 1159 249 1195 289
rect 1159 215 1210 249
rect 1244 215 1278 249
rect 1312 215 1346 249
rect 1380 215 1414 249
rect 1448 215 1464 249
rect 693 161 695 169
rect 36 135 695 161
rect 729 135 731 169
rect 1498 161 1547 293
rect 36 127 731 135
rect 36 101 88 127
rect 36 67 52 101
rect 86 67 88 101
rect 222 123 731 127
rect 765 123 781 157
rect 815 123 1099 157
rect 222 101 268 123
rect 36 51 88 67
rect 122 59 138 93
rect 172 59 188 93
rect 122 17 188 59
rect 222 67 224 101
rect 258 67 268 101
rect 403 101 448 123
rect 222 51 268 67
rect 302 55 318 89
rect 352 55 368 89
rect 302 17 368 55
rect 437 67 448 101
rect 693 101 731 123
rect 403 51 448 67
rect 484 55 500 89
rect 534 55 604 89
rect 638 55 659 89
rect 484 17 659 55
rect 693 67 695 101
rect 729 89 731 101
rect 1062 101 1099 123
rect 1233 127 1547 161
rect 729 67 866 89
rect 693 55 866 67
rect 900 55 917 89
rect 693 51 917 55
rect 961 55 978 89
rect 1012 55 1028 89
rect 961 17 1028 55
rect 1062 67 1063 101
rect 1097 67 1099 101
rect 1062 51 1099 67
rect 1133 89 1199 103
rect 1133 55 1149 89
rect 1183 55 1199 89
rect 1133 17 1199 55
rect 1233 101 1271 127
rect 1233 67 1235 101
rect 1269 67 1271 101
rect 1405 101 1443 127
rect 1233 51 1271 67
rect 1305 55 1321 89
rect 1355 55 1371 89
rect 1305 17 1371 55
rect 1405 67 1407 101
rect 1441 67 1443 101
rect 1405 51 1443 67
rect 1477 59 1493 93
rect 1527 59 1543 93
rect 1477 17 1543 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
<< metal1 >>
rect 0 561 1564 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 0 496 1564 527
rect 0 17 1564 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
rect 0 -48 1564 -17
<< labels >>
flabel locali s 305 221 339 255 0 FreeSans 400 0 0 0 C1
port 4 nsew signal input
flabel locali s 583 221 617 255 0 FreeSans 400 0 0 0 B1
port 3 nsew signal input
flabel locali s 859 221 893 255 0 FreeSans 400 0 0 0 A1
port 1 nsew signal input
flabel locali s 1045 221 1079 255 0 FreeSans 400 0 0 0 A2
port 2 nsew signal input
flabel locali s 1505 153 1539 187 0 FreeSans 400 0 0 0 X
port 10 nsew signal output
flabel locali s 29 221 63 255 0 FreeSans 400 0 0 0 D1
port 5 nsew signal input
flabel locali s 29 289 63 323 0 FreeSans 400 0 0 0 D1
port 5 nsew signal input
flabel locali s 213 221 247 255 0 FreeSans 400 0 0 0 C1
port 4 nsew signal input
flabel locali s 397 221 431 255 0 FreeSans 400 0 0 0 C1
port 4 nsew signal input
flabel locali s 491 221 525 255 0 FreeSans 400 0 0 0 B1
port 3 nsew signal input
flabel locali s 767 221 801 255 0 FreeSans 400 0 0 0 A1
port 1 nsew signal input
flabel locali s 951 221 987 255 0 FreeSans 400 0 0 0 A2
port 2 nsew signal input
flabel locali s 1505 221 1539 255 0 FreeSans 400 0 0 0 X
port 10 nsew signal output
flabel locali s 1505 289 1539 323 0 FreeSans 400 0 0 0 X
port 10 nsew signal output
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 a2111o_4
rlabel metal1 s 0 -48 1564 48 1 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1564 592 1 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1564 544
string GDS_END 3783064
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3770710
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 39.100 0.000 
<< end >>
