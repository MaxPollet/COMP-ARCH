magic
tech sky130A
magscale 1 2
timestamp 1681267127
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_0
timestamp 1681267127
transform 1 0 -50 0 1 13
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_1
timestamp 1681267127
transform 1 0 -50 0 1 -243
box 0 0 1 1
<< properties >>
string GDS_END 31311484
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 31310700
<< end >>
