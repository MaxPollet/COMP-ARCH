magic
tech sky130A
magscale 1 2
timestamp 1681267127
<< nwell >>
rect 0 0 524 1214
<< pmos >>
rect 204 102 234 1112
rect 290 102 320 1112
<< pdiff >>
rect 148 1100 204 1112
rect 148 1066 159 1100
rect 193 1066 204 1100
rect 148 1032 204 1066
rect 148 998 159 1032
rect 193 998 204 1032
rect 148 964 204 998
rect 148 930 159 964
rect 193 930 204 964
rect 148 896 204 930
rect 148 862 159 896
rect 193 862 204 896
rect 148 828 204 862
rect 148 794 159 828
rect 193 794 204 828
rect 148 760 204 794
rect 148 726 159 760
rect 193 726 204 760
rect 148 692 204 726
rect 148 658 159 692
rect 193 658 204 692
rect 148 624 204 658
rect 148 590 159 624
rect 193 590 204 624
rect 148 556 204 590
rect 148 522 159 556
rect 193 522 204 556
rect 148 488 204 522
rect 148 454 159 488
rect 193 454 204 488
rect 148 420 204 454
rect 148 386 159 420
rect 193 386 204 420
rect 148 352 204 386
rect 148 318 159 352
rect 193 318 204 352
rect 148 284 204 318
rect 148 250 159 284
rect 193 250 204 284
rect 148 216 204 250
rect 148 182 159 216
rect 193 182 204 216
rect 148 148 204 182
rect 148 114 159 148
rect 193 114 204 148
rect 148 102 204 114
rect 234 1100 290 1112
rect 234 1066 245 1100
rect 279 1066 290 1100
rect 234 1032 290 1066
rect 234 998 245 1032
rect 279 998 290 1032
rect 234 964 290 998
rect 234 930 245 964
rect 279 930 290 964
rect 234 896 290 930
rect 234 862 245 896
rect 279 862 290 896
rect 234 828 290 862
rect 234 794 245 828
rect 279 794 290 828
rect 234 760 290 794
rect 234 726 245 760
rect 279 726 290 760
rect 234 692 290 726
rect 234 658 245 692
rect 279 658 290 692
rect 234 624 290 658
rect 234 590 245 624
rect 279 590 290 624
rect 234 556 290 590
rect 234 522 245 556
rect 279 522 290 556
rect 234 488 290 522
rect 234 454 245 488
rect 279 454 290 488
rect 234 420 290 454
rect 234 386 245 420
rect 279 386 290 420
rect 234 352 290 386
rect 234 318 245 352
rect 279 318 290 352
rect 234 284 290 318
rect 234 250 245 284
rect 279 250 290 284
rect 234 216 290 250
rect 234 182 245 216
rect 279 182 290 216
rect 234 148 290 182
rect 234 114 245 148
rect 279 114 290 148
rect 234 102 290 114
rect 320 1100 376 1112
rect 320 1066 331 1100
rect 365 1066 376 1100
rect 320 1032 376 1066
rect 320 998 331 1032
rect 365 998 376 1032
rect 320 964 376 998
rect 320 930 331 964
rect 365 930 376 964
rect 320 896 376 930
rect 320 862 331 896
rect 365 862 376 896
rect 320 828 376 862
rect 320 794 331 828
rect 365 794 376 828
rect 320 760 376 794
rect 320 726 331 760
rect 365 726 376 760
rect 320 692 376 726
rect 320 658 331 692
rect 365 658 376 692
rect 320 624 376 658
rect 320 590 331 624
rect 365 590 376 624
rect 320 556 376 590
rect 320 522 331 556
rect 365 522 376 556
rect 320 488 376 522
rect 320 454 331 488
rect 365 454 376 488
rect 320 420 376 454
rect 320 386 331 420
rect 365 386 376 420
rect 320 352 376 386
rect 320 318 331 352
rect 365 318 376 352
rect 320 284 376 318
rect 320 250 331 284
rect 365 250 376 284
rect 320 216 376 250
rect 320 182 331 216
rect 365 182 376 216
rect 320 148 376 182
rect 320 114 331 148
rect 365 114 376 148
rect 320 102 376 114
<< pdiffc >>
rect 159 1066 193 1100
rect 159 998 193 1032
rect 159 930 193 964
rect 159 862 193 896
rect 159 794 193 828
rect 159 726 193 760
rect 159 658 193 692
rect 159 590 193 624
rect 159 522 193 556
rect 159 454 193 488
rect 159 386 193 420
rect 159 318 193 352
rect 159 250 193 284
rect 159 182 193 216
rect 159 114 193 148
rect 245 1066 279 1100
rect 245 998 279 1032
rect 245 930 279 964
rect 245 862 279 896
rect 245 794 279 828
rect 245 726 279 760
rect 245 658 279 692
rect 245 590 279 624
rect 245 522 279 556
rect 245 454 279 488
rect 245 386 279 420
rect 245 318 279 352
rect 245 250 279 284
rect 245 182 279 216
rect 245 114 279 148
rect 331 1066 365 1100
rect 331 998 365 1032
rect 331 930 365 964
rect 331 862 365 896
rect 331 794 365 828
rect 331 726 365 760
rect 331 658 365 692
rect 331 590 365 624
rect 331 522 365 556
rect 331 454 365 488
rect 331 386 365 420
rect 331 318 365 352
rect 331 250 365 284
rect 331 182 365 216
rect 331 114 365 148
<< nsubdiff >>
rect 36 1066 94 1112
rect 36 1032 48 1066
rect 82 1032 94 1066
rect 36 998 94 1032
rect 36 964 48 998
rect 82 964 94 998
rect 36 930 94 964
rect 36 896 48 930
rect 82 896 94 930
rect 36 862 94 896
rect 36 828 48 862
rect 82 828 94 862
rect 36 794 94 828
rect 36 760 48 794
rect 82 760 94 794
rect 36 726 94 760
rect 36 692 48 726
rect 82 692 94 726
rect 36 658 94 692
rect 36 624 48 658
rect 82 624 94 658
rect 36 590 94 624
rect 36 556 48 590
rect 82 556 94 590
rect 36 522 94 556
rect 36 488 48 522
rect 82 488 94 522
rect 36 454 94 488
rect 36 420 48 454
rect 82 420 94 454
rect 36 386 94 420
rect 36 352 48 386
rect 82 352 94 386
rect 36 318 94 352
rect 36 284 48 318
rect 82 284 94 318
rect 36 250 94 284
rect 36 216 48 250
rect 82 216 94 250
rect 36 182 94 216
rect 36 148 48 182
rect 82 148 94 182
rect 36 102 94 148
rect 430 1066 488 1112
rect 430 1032 442 1066
rect 476 1032 488 1066
rect 430 998 488 1032
rect 430 964 442 998
rect 476 964 488 998
rect 430 930 488 964
rect 430 896 442 930
rect 476 896 488 930
rect 430 862 488 896
rect 430 828 442 862
rect 476 828 488 862
rect 430 794 488 828
rect 430 760 442 794
rect 476 760 488 794
rect 430 726 488 760
rect 430 692 442 726
rect 476 692 488 726
rect 430 658 488 692
rect 430 624 442 658
rect 476 624 488 658
rect 430 590 488 624
rect 430 556 442 590
rect 476 556 488 590
rect 430 522 488 556
rect 430 488 442 522
rect 476 488 488 522
rect 430 454 488 488
rect 430 420 442 454
rect 476 420 488 454
rect 430 386 488 420
rect 430 352 442 386
rect 476 352 488 386
rect 430 318 488 352
rect 430 284 442 318
rect 476 284 488 318
rect 430 250 488 284
rect 430 216 442 250
rect 476 216 488 250
rect 430 182 488 216
rect 430 148 442 182
rect 476 148 488 182
rect 430 102 488 148
<< nsubdiffcont >>
rect 48 1032 82 1066
rect 48 964 82 998
rect 48 896 82 930
rect 48 828 82 862
rect 48 760 82 794
rect 48 692 82 726
rect 48 624 82 658
rect 48 556 82 590
rect 48 488 82 522
rect 48 420 82 454
rect 48 352 82 386
rect 48 284 82 318
rect 48 216 82 250
rect 48 148 82 182
rect 442 1032 476 1066
rect 442 964 476 998
rect 442 896 476 930
rect 442 828 476 862
rect 442 760 476 794
rect 442 692 476 726
rect 442 624 476 658
rect 442 556 476 590
rect 442 488 476 522
rect 442 420 476 454
rect 442 352 476 386
rect 442 284 476 318
rect 442 216 476 250
rect 442 148 476 182
<< poly >>
rect 161 1194 363 1214
rect 161 1160 177 1194
rect 211 1160 245 1194
rect 279 1160 313 1194
rect 347 1160 363 1194
rect 161 1144 363 1160
rect 161 54 363 70
rect 161 20 177 54
rect 211 20 245 54
rect 279 20 313 54
rect 347 20 363 54
rect 161 0 363 20
<< polycont >>
rect 177 1160 211 1194
rect 245 1160 279 1194
rect 313 1160 347 1194
rect 177 20 211 54
rect 245 20 279 54
rect 313 20 347 54
<< locali >>
rect 161 1160 173 1194
rect 211 1160 245 1194
rect 279 1160 313 1194
rect 351 1160 363 1194
rect 159 1100 193 1116
rect 48 1020 82 1032
rect 48 948 82 964
rect 48 876 82 896
rect 48 804 82 828
rect 48 732 82 760
rect 48 660 82 692
rect 48 590 82 624
rect 48 522 82 554
rect 48 454 82 482
rect 48 386 82 410
rect 48 318 82 338
rect 48 250 82 266
rect 48 182 82 194
rect 159 1032 193 1058
rect 159 964 193 986
rect 159 896 193 914
rect 159 828 193 842
rect 159 760 193 770
rect 159 692 193 698
rect 159 624 193 626
rect 159 588 193 590
rect 159 516 193 522
rect 159 444 193 454
rect 159 372 193 386
rect 159 300 193 318
rect 159 228 193 250
rect 159 156 193 182
rect 159 98 193 114
rect 245 1100 279 1116
rect 245 1032 279 1058
rect 245 964 279 986
rect 245 896 279 914
rect 245 828 279 842
rect 245 760 279 770
rect 245 692 279 698
rect 245 624 279 626
rect 245 588 279 590
rect 245 516 279 522
rect 245 444 279 454
rect 245 372 279 386
rect 245 300 279 318
rect 245 228 279 250
rect 245 156 279 182
rect 245 98 279 114
rect 331 1100 365 1116
rect 331 1032 365 1058
rect 331 964 365 986
rect 331 896 365 914
rect 331 828 365 842
rect 331 760 365 770
rect 331 692 365 698
rect 331 624 365 626
rect 331 588 365 590
rect 331 516 365 522
rect 331 444 365 454
rect 331 372 365 386
rect 331 300 365 318
rect 331 228 365 250
rect 331 156 365 182
rect 442 1020 476 1032
rect 442 948 476 964
rect 442 876 476 896
rect 442 804 476 828
rect 442 732 476 760
rect 442 660 476 692
rect 442 590 476 624
rect 442 522 476 554
rect 442 454 476 482
rect 442 386 476 410
rect 442 318 476 338
rect 442 250 476 266
rect 442 182 476 194
rect 331 98 365 114
rect 161 20 173 54
rect 211 20 245 54
rect 279 20 313 54
rect 351 20 363 54
<< viali >>
rect 173 1160 177 1194
rect 177 1160 207 1194
rect 245 1160 279 1194
rect 317 1160 347 1194
rect 347 1160 351 1194
rect 48 1066 82 1092
rect 48 1058 82 1066
rect 48 998 82 1020
rect 48 986 82 998
rect 48 930 82 948
rect 48 914 82 930
rect 48 862 82 876
rect 48 842 82 862
rect 48 794 82 804
rect 48 770 82 794
rect 48 726 82 732
rect 48 698 82 726
rect 48 658 82 660
rect 48 626 82 658
rect 48 556 82 588
rect 48 554 82 556
rect 48 488 82 516
rect 48 482 82 488
rect 48 420 82 444
rect 48 410 82 420
rect 48 352 82 372
rect 48 338 82 352
rect 48 284 82 300
rect 48 266 82 284
rect 48 216 82 228
rect 48 194 82 216
rect 48 148 82 156
rect 48 122 82 148
rect 159 1066 193 1092
rect 159 1058 193 1066
rect 159 998 193 1020
rect 159 986 193 998
rect 159 930 193 948
rect 159 914 193 930
rect 159 862 193 876
rect 159 842 193 862
rect 159 794 193 804
rect 159 770 193 794
rect 159 726 193 732
rect 159 698 193 726
rect 159 658 193 660
rect 159 626 193 658
rect 159 556 193 588
rect 159 554 193 556
rect 159 488 193 516
rect 159 482 193 488
rect 159 420 193 444
rect 159 410 193 420
rect 159 352 193 372
rect 159 338 193 352
rect 159 284 193 300
rect 159 266 193 284
rect 159 216 193 228
rect 159 194 193 216
rect 159 148 193 156
rect 159 122 193 148
rect 245 1066 279 1092
rect 245 1058 279 1066
rect 245 998 279 1020
rect 245 986 279 998
rect 245 930 279 948
rect 245 914 279 930
rect 245 862 279 876
rect 245 842 279 862
rect 245 794 279 804
rect 245 770 279 794
rect 245 726 279 732
rect 245 698 279 726
rect 245 658 279 660
rect 245 626 279 658
rect 245 556 279 588
rect 245 554 279 556
rect 245 488 279 516
rect 245 482 279 488
rect 245 420 279 444
rect 245 410 279 420
rect 245 352 279 372
rect 245 338 279 352
rect 245 284 279 300
rect 245 266 279 284
rect 245 216 279 228
rect 245 194 279 216
rect 245 148 279 156
rect 245 122 279 148
rect 331 1066 365 1092
rect 331 1058 365 1066
rect 331 998 365 1020
rect 331 986 365 998
rect 331 930 365 948
rect 331 914 365 930
rect 331 862 365 876
rect 331 842 365 862
rect 331 794 365 804
rect 331 770 365 794
rect 331 726 365 732
rect 331 698 365 726
rect 331 658 365 660
rect 331 626 365 658
rect 331 556 365 588
rect 331 554 365 556
rect 331 488 365 516
rect 331 482 365 488
rect 331 420 365 444
rect 331 410 365 420
rect 331 352 365 372
rect 331 338 365 352
rect 331 284 365 300
rect 331 266 365 284
rect 331 216 365 228
rect 331 194 365 216
rect 331 148 365 156
rect 331 122 365 148
rect 442 1066 476 1092
rect 442 1058 476 1066
rect 442 998 476 1020
rect 442 986 476 998
rect 442 930 476 948
rect 442 914 476 930
rect 442 862 476 876
rect 442 842 476 862
rect 442 794 476 804
rect 442 770 476 794
rect 442 726 476 732
rect 442 698 476 726
rect 442 658 476 660
rect 442 626 476 658
rect 442 556 476 588
rect 442 554 476 556
rect 442 488 476 516
rect 442 482 476 488
rect 442 420 476 444
rect 442 410 476 420
rect 442 352 476 372
rect 442 338 476 352
rect 442 284 476 300
rect 442 266 476 284
rect 442 216 476 228
rect 442 194 476 216
rect 442 148 476 156
rect 442 122 476 148
rect 173 20 177 54
rect 177 20 207 54
rect 245 20 279 54
rect 317 20 347 54
rect 347 20 351 54
<< metal1 >>
rect 161 1194 363 1214
rect 161 1160 173 1194
rect 207 1160 245 1194
rect 279 1160 317 1194
rect 351 1160 363 1194
rect 161 1148 363 1160
rect 36 1092 94 1104
rect 36 1058 48 1092
rect 82 1058 94 1092
rect 36 1020 94 1058
rect 36 986 48 1020
rect 82 986 94 1020
rect 36 948 94 986
rect 36 914 48 948
rect 82 914 94 948
rect 36 876 94 914
rect 36 842 48 876
rect 82 842 94 876
rect 36 804 94 842
rect 36 770 48 804
rect 82 770 94 804
rect 36 732 94 770
rect 36 698 48 732
rect 82 698 94 732
rect 36 660 94 698
rect 36 626 48 660
rect 82 626 94 660
rect 36 588 94 626
rect 36 554 48 588
rect 82 554 94 588
rect 36 516 94 554
rect 36 482 48 516
rect 82 482 94 516
rect 36 444 94 482
rect 36 410 48 444
rect 82 410 94 444
rect 36 372 94 410
rect 36 338 48 372
rect 82 338 94 372
rect 36 300 94 338
rect 36 266 48 300
rect 82 266 94 300
rect 36 228 94 266
rect 36 194 48 228
rect 82 194 94 228
rect 36 156 94 194
rect 36 122 48 156
rect 82 122 94 156
rect 36 110 94 122
rect 150 1092 202 1104
rect 150 1058 159 1092
rect 193 1058 202 1092
rect 150 1020 202 1058
rect 150 986 159 1020
rect 193 986 202 1020
rect 150 948 202 986
rect 150 914 159 948
rect 193 914 202 948
rect 150 876 202 914
rect 150 842 159 876
rect 193 842 202 876
rect 150 804 202 842
rect 150 770 159 804
rect 193 770 202 804
rect 150 732 202 770
rect 150 698 159 732
rect 193 698 202 732
rect 150 660 202 698
rect 150 626 159 660
rect 193 626 202 660
rect 150 588 202 626
rect 150 554 159 588
rect 193 554 202 588
rect 150 552 202 554
rect 150 488 159 500
rect 193 488 202 500
rect 150 424 159 436
rect 193 424 202 436
rect 150 360 159 372
rect 193 360 202 372
rect 150 300 202 308
rect 150 296 159 300
rect 193 296 202 300
rect 150 232 202 244
rect 150 168 202 180
rect 150 110 202 116
rect 236 1098 288 1104
rect 236 1034 288 1046
rect 236 970 288 982
rect 236 914 245 918
rect 279 914 288 918
rect 236 906 288 914
rect 236 842 245 854
rect 279 842 288 854
rect 236 778 245 790
rect 279 778 288 790
rect 236 714 245 726
rect 279 714 288 726
rect 236 660 288 662
rect 236 626 245 660
rect 279 626 288 660
rect 236 588 288 626
rect 236 554 245 588
rect 279 554 288 588
rect 236 516 288 554
rect 236 482 245 516
rect 279 482 288 516
rect 236 444 288 482
rect 236 410 245 444
rect 279 410 288 444
rect 236 372 288 410
rect 236 338 245 372
rect 279 338 288 372
rect 236 300 288 338
rect 236 266 245 300
rect 279 266 288 300
rect 236 228 288 266
rect 236 194 245 228
rect 279 194 288 228
rect 236 156 288 194
rect 236 122 245 156
rect 279 122 288 156
rect 236 110 288 122
rect 322 1092 374 1104
rect 322 1058 331 1092
rect 365 1058 374 1092
rect 322 1020 374 1058
rect 322 986 331 1020
rect 365 986 374 1020
rect 322 948 374 986
rect 322 914 331 948
rect 365 914 374 948
rect 322 876 374 914
rect 322 842 331 876
rect 365 842 374 876
rect 322 804 374 842
rect 322 770 331 804
rect 365 770 374 804
rect 322 732 374 770
rect 322 698 331 732
rect 365 698 374 732
rect 322 660 374 698
rect 322 626 331 660
rect 365 626 374 660
rect 322 588 374 626
rect 322 554 331 588
rect 365 554 374 588
rect 322 552 374 554
rect 322 488 331 500
rect 365 488 374 500
rect 322 424 331 436
rect 365 424 374 436
rect 322 360 331 372
rect 365 360 374 372
rect 322 300 374 308
rect 322 296 331 300
rect 365 296 374 300
rect 322 232 374 244
rect 322 168 374 180
rect 322 110 374 116
rect 430 1092 488 1104
rect 430 1058 442 1092
rect 476 1058 488 1092
rect 430 1020 488 1058
rect 430 986 442 1020
rect 476 986 488 1020
rect 430 948 488 986
rect 430 914 442 948
rect 476 914 488 948
rect 430 876 488 914
rect 430 842 442 876
rect 476 842 488 876
rect 430 804 488 842
rect 430 770 442 804
rect 476 770 488 804
rect 430 732 488 770
rect 430 698 442 732
rect 476 698 488 732
rect 430 660 488 698
rect 430 626 442 660
rect 476 626 488 660
rect 430 588 488 626
rect 430 554 442 588
rect 476 554 488 588
rect 430 516 488 554
rect 430 482 442 516
rect 476 482 488 516
rect 430 444 488 482
rect 430 410 442 444
rect 476 410 488 444
rect 430 372 488 410
rect 430 338 442 372
rect 476 338 488 372
rect 430 300 488 338
rect 430 266 442 300
rect 476 266 488 300
rect 430 228 488 266
rect 430 194 442 228
rect 476 194 488 228
rect 430 156 488 194
rect 430 122 442 156
rect 476 122 488 156
rect 430 110 488 122
rect 161 54 363 66
rect 161 20 173 54
rect 207 20 245 54
rect 279 20 317 54
rect 351 20 363 54
rect 161 0 363 20
<< via1 >>
rect 150 516 202 552
rect 150 500 159 516
rect 159 500 193 516
rect 193 500 202 516
rect 150 482 159 488
rect 159 482 193 488
rect 193 482 202 488
rect 150 444 202 482
rect 150 436 159 444
rect 159 436 193 444
rect 193 436 202 444
rect 150 410 159 424
rect 159 410 193 424
rect 193 410 202 424
rect 150 372 202 410
rect 150 338 159 360
rect 159 338 193 360
rect 193 338 202 360
rect 150 308 202 338
rect 150 266 159 296
rect 159 266 193 296
rect 193 266 202 296
rect 150 244 202 266
rect 150 228 202 232
rect 150 194 159 228
rect 159 194 193 228
rect 193 194 202 228
rect 150 180 202 194
rect 150 156 202 168
rect 150 122 159 156
rect 159 122 193 156
rect 193 122 202 156
rect 150 116 202 122
rect 236 1092 288 1098
rect 236 1058 245 1092
rect 245 1058 279 1092
rect 279 1058 288 1092
rect 236 1046 288 1058
rect 236 1020 288 1034
rect 236 986 245 1020
rect 245 986 279 1020
rect 279 986 288 1020
rect 236 982 288 986
rect 236 948 288 970
rect 236 918 245 948
rect 245 918 279 948
rect 279 918 288 948
rect 236 876 288 906
rect 236 854 245 876
rect 245 854 279 876
rect 279 854 288 876
rect 236 804 288 842
rect 236 790 245 804
rect 245 790 279 804
rect 279 790 288 804
rect 236 770 245 778
rect 245 770 279 778
rect 279 770 288 778
rect 236 732 288 770
rect 236 726 245 732
rect 245 726 279 732
rect 279 726 288 732
rect 236 698 245 714
rect 245 698 279 714
rect 279 698 288 714
rect 236 662 288 698
rect 322 516 374 552
rect 322 500 331 516
rect 331 500 365 516
rect 365 500 374 516
rect 322 482 331 488
rect 331 482 365 488
rect 365 482 374 488
rect 322 444 374 482
rect 322 436 331 444
rect 331 436 365 444
rect 365 436 374 444
rect 322 410 331 424
rect 331 410 365 424
rect 365 410 374 424
rect 322 372 374 410
rect 322 338 331 360
rect 331 338 365 360
rect 365 338 374 360
rect 322 308 374 338
rect 322 266 331 296
rect 331 266 365 296
rect 365 266 374 296
rect 322 244 374 266
rect 322 228 374 232
rect 322 194 331 228
rect 331 194 365 228
rect 365 194 374 228
rect 322 180 374 194
rect 322 156 374 168
rect 322 122 331 156
rect 331 122 365 156
rect 365 122 374 156
rect 322 116 374 122
<< metal2 >>
rect 10 1098 514 1104
rect 10 1046 236 1098
rect 288 1046 514 1098
rect 10 1034 514 1046
rect 10 982 236 1034
rect 288 982 514 1034
rect 10 970 514 982
rect 10 918 236 970
rect 288 918 514 970
rect 10 906 514 918
rect 10 854 236 906
rect 288 854 514 906
rect 10 842 514 854
rect 10 790 236 842
rect 288 790 514 842
rect 10 778 514 790
rect 10 726 236 778
rect 288 726 514 778
rect 10 714 514 726
rect 10 662 236 714
rect 288 662 514 714
rect 10 632 514 662
rect 10 552 514 582
rect 10 500 150 552
rect 202 500 322 552
rect 374 500 514 552
rect 10 488 514 500
rect 10 436 150 488
rect 202 436 322 488
rect 374 436 514 488
rect 10 424 514 436
rect 10 372 150 424
rect 202 372 322 424
rect 374 372 514 424
rect 10 360 514 372
rect 10 308 150 360
rect 202 308 322 360
rect 374 308 514 360
rect 10 296 514 308
rect 10 244 150 296
rect 202 244 322 296
rect 374 244 514 296
rect 10 232 514 244
rect 10 180 150 232
rect 202 180 322 232
rect 374 180 514 232
rect 10 168 514 180
rect 10 116 150 168
rect 202 116 322 168
rect 374 116 514 168
rect 10 110 514 116
<< labels >>
flabel metal2 s 10 632 30 1104 7 FreeSans 300 180 0 0 DRAIN
port 2 nsew
flabel metal2 s 10 110 30 582 7 FreeSans 300 180 0 0 SOURCE
port 3 nsew
flabel metal1 s 430 110 488 126 3 FreeSans 300 90 0 0 BULK
port 4 nsew
flabel metal1 s 161 1148 363 1214 0 FreeSans 300 0 0 0 GATE
port 5 nsew
flabel metal1 s 161 0 363 66 0 FreeSans 300 0 0 0 GATE
port 5 nsew
flabel metal1 s 36 110 94 126 3 FreeSans 300 90 0 0 BULK
port 4 nsew
<< properties >>
string GDS_END 9362650
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 9347190
<< end >>
