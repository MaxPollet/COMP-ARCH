magic
tech sky130A
magscale 1 2
timestamp 1681267127
<< nwell >>
rect -66 377 930 897
<< pwell >>
rect 20 43 856 283
rect -26 -43 890 43
<< mvnmos >>
rect 103 107 203 257
rect 375 107 475 257
rect 531 107 631 257
rect 673 107 773 257
<< mvpmos >>
rect 83 443 183 743
rect 369 443 469 743
rect 525 443 625 743
rect 681 443 781 743
<< mvndiff >>
rect 46 249 103 257
rect 46 215 58 249
rect 92 215 103 249
rect 46 149 103 215
rect 46 115 58 149
rect 92 115 103 149
rect 46 107 103 115
rect 203 249 375 257
rect 203 215 214 249
rect 248 215 375 249
rect 203 149 375 215
rect 203 115 214 149
rect 248 115 375 149
rect 203 107 375 115
rect 475 249 531 257
rect 475 215 486 249
rect 520 215 531 249
rect 475 149 531 215
rect 475 115 486 149
rect 520 115 531 149
rect 475 107 531 115
rect 631 107 673 257
rect 773 249 830 257
rect 773 215 784 249
rect 818 215 830 249
rect 773 149 830 215
rect 773 115 784 149
rect 818 115 830 149
rect 773 107 830 115
<< mvpdiff >>
rect 30 731 83 743
rect 30 697 38 731
rect 72 697 83 731
rect 30 651 83 697
rect 30 617 38 651
rect 72 617 83 651
rect 30 569 83 617
rect 30 535 38 569
rect 72 535 83 569
rect 30 489 83 535
rect 30 455 38 489
rect 72 455 83 489
rect 30 443 83 455
rect 183 735 240 743
rect 183 701 194 735
rect 228 701 240 735
rect 183 654 240 701
rect 183 620 194 654
rect 228 620 240 654
rect 183 571 240 620
rect 183 537 194 571
rect 228 537 240 571
rect 183 490 240 537
rect 183 456 194 490
rect 228 456 240 490
rect 183 443 240 456
rect 312 735 369 743
rect 312 701 324 735
rect 358 701 369 735
rect 312 652 369 701
rect 312 618 324 652
rect 358 618 369 652
rect 312 568 369 618
rect 312 534 324 568
rect 358 534 369 568
rect 312 485 369 534
rect 312 451 324 485
rect 358 451 369 485
rect 312 443 369 451
rect 469 735 525 743
rect 469 701 480 735
rect 514 701 525 735
rect 469 654 525 701
rect 469 620 480 654
rect 514 620 525 654
rect 469 571 525 620
rect 469 537 480 571
rect 514 537 525 571
rect 469 490 525 537
rect 469 456 480 490
rect 514 456 525 490
rect 469 443 525 456
rect 625 735 681 743
rect 625 701 636 735
rect 670 701 681 735
rect 625 647 681 701
rect 625 613 636 647
rect 670 613 681 647
rect 625 560 681 613
rect 625 526 636 560
rect 670 526 681 560
rect 625 443 681 526
rect 781 731 834 743
rect 781 697 792 731
rect 826 697 834 731
rect 781 651 834 697
rect 781 617 792 651
rect 826 617 834 651
rect 781 569 834 617
rect 781 535 792 569
rect 826 535 834 569
rect 781 489 834 535
rect 781 455 792 489
rect 826 455 834 489
rect 781 443 834 455
<< mvndiffc >>
rect 58 215 92 249
rect 58 115 92 149
rect 214 215 248 249
rect 214 115 248 149
rect 486 215 520 249
rect 486 115 520 149
rect 784 215 818 249
rect 784 115 818 149
<< mvpdiffc >>
rect 38 697 72 731
rect 38 617 72 651
rect 38 535 72 569
rect 38 455 72 489
rect 194 701 228 735
rect 194 620 228 654
rect 194 537 228 571
rect 194 456 228 490
rect 324 701 358 735
rect 324 618 358 652
rect 324 534 358 568
rect 324 451 358 485
rect 480 701 514 735
rect 480 620 514 654
rect 480 537 514 571
rect 480 456 514 490
rect 636 701 670 735
rect 636 613 670 647
rect 636 526 670 560
rect 792 697 826 731
rect 792 617 826 651
rect 792 535 826 569
rect 792 455 826 489
<< mvpsubdiff >>
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< mvnsubdiff >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 864 831
<< mvpsubdiffcont >>
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< mvnsubdiffcont >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
<< poly >>
rect 83 417 183 443
rect 83 395 203 417
rect 83 361 129 395
rect 163 361 203 395
rect 83 283 203 361
rect 369 383 469 443
rect 525 383 625 443
rect 681 417 781 443
rect 369 343 475 383
rect 369 309 389 343
rect 423 309 475 343
rect 369 283 475 309
rect 525 351 631 383
rect 525 317 577 351
rect 611 317 631 351
rect 525 283 631 317
rect 103 257 203 283
rect 375 257 475 283
rect 531 257 631 283
rect 673 351 843 417
rect 673 317 789 351
rect 823 317 843 351
rect 673 283 843 317
rect 673 257 773 283
<< polycont >>
rect 129 361 163 395
rect 389 309 423 343
rect 577 317 611 351
rect 789 317 823 351
<< locali >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 864 831
rect 22 731 72 747
rect 22 697 38 731
rect 22 651 72 697
rect 22 617 38 651
rect 22 569 72 617
rect 22 535 38 569
rect 22 489 72 535
rect 22 455 38 489
rect 108 735 288 751
rect 108 701 109 735
rect 143 701 181 735
rect 228 701 253 735
rect 287 701 288 735
rect 108 654 288 701
rect 108 620 194 654
rect 228 620 288 654
rect 108 571 288 620
rect 108 537 194 571
rect 228 537 288 571
rect 108 490 288 537
rect 108 456 194 490
rect 228 456 288 490
rect 324 735 374 751
rect 358 701 374 735
rect 324 652 374 701
rect 358 618 374 652
rect 324 568 374 618
rect 358 534 374 568
rect 324 485 374 534
rect 22 265 72 455
rect 358 451 374 485
rect 464 735 530 751
rect 464 701 480 735
rect 514 701 530 735
rect 464 654 530 701
rect 464 620 480 654
rect 514 620 530 654
rect 464 571 530 620
rect 464 537 480 571
rect 514 537 530 571
rect 464 490 530 537
rect 566 735 756 751
rect 566 701 572 735
rect 606 701 636 735
rect 678 701 716 735
rect 750 701 756 735
rect 566 647 756 701
rect 566 613 636 647
rect 670 613 756 647
rect 566 560 756 613
rect 566 526 636 560
rect 670 526 756 560
rect 792 731 842 747
rect 826 697 842 731
rect 792 651 842 697
rect 826 617 842 651
rect 792 569 842 617
rect 826 535 842 569
rect 792 490 842 535
rect 464 456 480 490
rect 514 489 842 490
rect 514 456 792 489
rect 324 420 374 451
rect 826 455 842 489
rect 792 439 842 455
rect 113 395 525 420
rect 113 361 129 395
rect 163 386 525 395
rect 163 361 179 386
rect 113 345 179 361
rect 217 343 455 350
rect 217 309 389 343
rect 423 309 455 343
rect 217 301 455 309
rect 491 265 525 386
rect 561 351 743 367
rect 561 317 577 351
rect 611 317 743 351
rect 561 301 743 317
rect 779 351 839 367
rect 779 317 789 351
rect 823 317 839 351
rect 779 301 839 317
rect 22 249 92 265
rect 22 215 58 249
rect 22 149 92 215
rect 22 115 58 149
rect 22 99 92 115
rect 128 249 450 265
rect 128 215 214 249
rect 248 215 450 249
rect 128 149 450 215
rect 128 115 214 149
rect 248 115 450 149
rect 128 113 450 115
rect 162 79 200 113
rect 234 79 272 113
rect 306 79 344 113
rect 378 79 416 113
rect 486 249 536 265
rect 520 215 536 249
rect 486 149 536 215
rect 520 115 536 149
rect 486 99 536 115
rect 572 249 834 265
rect 572 215 784 249
rect 818 215 834 249
rect 572 149 834 215
rect 572 115 784 149
rect 818 115 834 149
rect 572 113 834 115
rect 128 73 450 79
rect 572 79 578 113
rect 612 79 650 113
rect 684 79 722 113
rect 756 79 794 113
rect 828 79 834 113
rect 572 73 834 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 109 701 143 735
rect 181 701 194 735
rect 194 701 215 735
rect 253 701 287 735
rect 572 701 606 735
rect 644 701 670 735
rect 670 701 678 735
rect 716 701 750 735
rect 128 79 162 113
rect 200 79 234 113
rect 272 79 306 113
rect 344 79 378 113
rect 416 79 450 113
rect 578 79 612 113
rect 650 79 684 113
rect 722 79 756 113
rect 794 79 828 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 831 864 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 864 831
rect 0 791 864 797
rect 0 735 864 763
rect 0 701 109 735
rect 143 701 181 735
rect 215 701 253 735
rect 287 701 572 735
rect 606 701 644 735
rect 678 701 716 735
rect 750 701 864 735
rect 0 689 864 701
rect 0 113 864 125
rect 0 79 128 113
rect 162 79 200 113
rect 234 79 272 113
rect 306 79 344 113
rect 378 79 416 113
rect 450 79 578 113
rect 612 79 650 113
rect 684 79 722 113
rect 756 79 794 113
rect 828 79 864 113
rect 0 51 864 79
rect 0 17 864 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -23 864 -17
<< labels >>
rlabel comment s 0 0 0 0 4 a21o_1
flabel metal1 s 0 51 864 125 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel metal1 s 0 0 864 23 0 FreeSans 340 0 0 0 VNB
port 5 nsew ground bidirectional
flabel metal1 s 0 689 864 763 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 791 864 814 0 FreeSans 340 0 0 0 VPB
port 6 nsew power bidirectional
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 612 65 646 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 864 814
string GDS_END 760356
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 748722
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
<< end >>
