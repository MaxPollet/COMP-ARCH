magic
tech sky130A
magscale 1 2
timestamp 1681267127
<< nwell >>
rect -38 261 2062 582
<< pwell >>
rect 1 21 1991 203
rect 30 -17 64 21
<< scnmos >>
rect 83 47 113 177
rect 167 47 197 177
rect 253 47 283 177
rect 339 47 369 177
rect 441 47 471 177
rect 527 47 557 177
rect 613 47 643 177
rect 699 47 729 177
rect 807 47 837 177
rect 893 47 923 177
rect 979 47 1009 177
rect 1065 47 1095 177
rect 1261 47 1291 177
rect 1347 47 1377 177
rect 1433 47 1463 177
rect 1519 47 1549 177
rect 1624 47 1654 177
rect 1710 47 1740 177
rect 1796 47 1826 177
rect 1882 47 1912 177
<< scpmoshvt >>
rect 81 297 111 497
rect 167 297 197 497
rect 253 297 283 497
rect 339 297 369 497
rect 425 297 455 497
rect 511 297 541 497
rect 597 297 627 497
rect 683 297 713 497
rect 873 297 903 497
rect 959 297 989 497
rect 1045 297 1075 497
rect 1131 297 1161 497
rect 1219 297 1249 497
rect 1305 297 1335 497
rect 1391 297 1421 497
rect 1481 297 1511 497
rect 1591 297 1621 497
rect 1677 297 1707 497
rect 1781 297 1811 497
rect 1867 297 1897 497
<< ndiff >>
rect 27 89 83 177
rect 27 55 39 89
rect 73 55 83 89
rect 27 47 83 55
rect 113 141 167 177
rect 113 107 123 141
rect 157 107 167 141
rect 113 47 167 107
rect 197 89 253 177
rect 197 55 208 89
rect 242 55 253 89
rect 197 47 253 55
rect 283 141 339 177
rect 283 107 294 141
rect 328 107 339 141
rect 283 47 339 107
rect 369 89 441 177
rect 369 55 396 89
rect 430 55 441 89
rect 369 47 441 55
rect 471 141 527 177
rect 471 107 482 141
rect 516 107 527 141
rect 471 47 527 107
rect 557 89 613 177
rect 557 55 568 89
rect 602 55 613 89
rect 557 47 613 55
rect 643 141 699 177
rect 643 107 654 141
rect 688 107 699 141
rect 643 47 699 107
rect 729 89 807 177
rect 729 55 752 89
rect 786 55 807 89
rect 729 47 807 55
rect 837 141 893 177
rect 837 107 848 141
rect 882 107 893 141
rect 837 47 893 107
rect 923 89 979 177
rect 923 55 934 89
rect 968 55 979 89
rect 923 47 979 55
rect 1009 141 1065 177
rect 1009 107 1020 141
rect 1054 107 1065 141
rect 1009 47 1065 107
rect 1095 89 1151 177
rect 1095 55 1105 89
rect 1139 55 1151 89
rect 1095 47 1151 55
rect 1205 89 1261 177
rect 1205 55 1217 89
rect 1251 55 1261 89
rect 1205 47 1261 55
rect 1291 157 1347 177
rect 1291 123 1302 157
rect 1336 123 1347 157
rect 1291 47 1347 123
rect 1377 89 1433 177
rect 1377 55 1388 89
rect 1422 55 1433 89
rect 1377 47 1433 55
rect 1463 157 1519 177
rect 1463 123 1474 157
rect 1508 123 1519 157
rect 1463 47 1519 123
rect 1549 119 1624 177
rect 1549 85 1578 119
rect 1612 85 1624 119
rect 1549 47 1624 85
rect 1654 89 1710 177
rect 1654 55 1665 89
rect 1699 55 1710 89
rect 1654 47 1710 55
rect 1740 119 1796 177
rect 1740 85 1751 119
rect 1785 85 1796 119
rect 1740 47 1796 85
rect 1826 89 1882 177
rect 1826 55 1837 89
rect 1871 55 1882 89
rect 1826 47 1882 55
rect 1912 119 1965 177
rect 1912 85 1923 119
rect 1957 85 1965 119
rect 1912 47 1965 85
<< pdiff >>
rect 28 485 81 497
rect 28 451 36 485
rect 70 451 81 485
rect 28 417 81 451
rect 28 383 36 417
rect 70 383 81 417
rect 28 297 81 383
rect 111 413 167 497
rect 111 379 122 413
rect 156 379 167 413
rect 111 345 167 379
rect 111 311 122 345
rect 156 311 167 345
rect 111 297 167 311
rect 197 489 253 497
rect 197 455 208 489
rect 242 455 253 489
rect 197 421 253 455
rect 197 387 208 421
rect 242 387 253 421
rect 197 297 253 387
rect 283 417 339 497
rect 283 383 294 417
rect 328 383 339 417
rect 283 348 339 383
rect 283 314 294 348
rect 328 314 339 348
rect 283 297 339 314
rect 369 489 425 497
rect 369 455 380 489
rect 414 455 425 489
rect 369 421 425 455
rect 369 387 380 421
rect 414 387 425 421
rect 369 297 425 387
rect 455 417 511 497
rect 455 383 466 417
rect 500 383 511 417
rect 455 349 511 383
rect 455 315 466 349
rect 500 315 511 349
rect 455 297 511 315
rect 541 489 597 497
rect 541 455 552 489
rect 586 455 597 489
rect 541 421 597 455
rect 541 387 552 421
rect 586 387 597 421
rect 541 297 597 387
rect 627 417 683 497
rect 627 383 638 417
rect 672 383 683 417
rect 627 348 683 383
rect 627 314 638 348
rect 672 314 683 348
rect 627 297 683 314
rect 713 485 765 497
rect 713 451 723 485
rect 757 451 765 485
rect 713 417 765 451
rect 713 383 723 417
rect 757 383 765 417
rect 713 297 765 383
rect 821 485 873 497
rect 821 451 829 485
rect 863 451 873 485
rect 821 417 873 451
rect 821 383 829 417
rect 863 383 873 417
rect 821 297 873 383
rect 903 417 959 497
rect 903 383 914 417
rect 948 383 959 417
rect 903 348 959 383
rect 903 314 914 348
rect 948 314 959 348
rect 903 297 959 314
rect 989 489 1045 497
rect 989 455 1000 489
rect 1034 455 1045 489
rect 989 421 1045 455
rect 989 387 1000 421
rect 1034 387 1045 421
rect 989 297 1045 387
rect 1075 417 1131 497
rect 1075 383 1086 417
rect 1120 383 1131 417
rect 1075 348 1131 383
rect 1075 314 1086 348
rect 1120 314 1131 348
rect 1075 297 1131 314
rect 1161 473 1219 497
rect 1161 439 1174 473
rect 1208 439 1219 473
rect 1161 343 1219 439
rect 1161 309 1174 343
rect 1208 309 1219 343
rect 1161 297 1219 309
rect 1249 489 1305 497
rect 1249 455 1260 489
rect 1294 455 1305 489
rect 1249 395 1305 455
rect 1249 361 1260 395
rect 1294 361 1305 395
rect 1249 297 1305 361
rect 1335 437 1391 497
rect 1335 403 1346 437
rect 1380 403 1391 437
rect 1335 343 1391 403
rect 1335 309 1346 343
rect 1380 309 1391 343
rect 1335 297 1391 309
rect 1421 489 1481 497
rect 1421 455 1432 489
rect 1466 455 1481 489
rect 1421 395 1481 455
rect 1421 361 1432 395
rect 1466 361 1481 395
rect 1421 297 1481 361
rect 1511 442 1591 497
rect 1511 408 1532 442
rect 1566 408 1591 442
rect 1511 343 1591 408
rect 1511 309 1522 343
rect 1556 309 1591 343
rect 1511 297 1591 309
rect 1621 485 1677 497
rect 1621 451 1632 485
rect 1666 451 1677 485
rect 1621 413 1677 451
rect 1621 379 1632 413
rect 1666 379 1677 413
rect 1621 297 1677 379
rect 1707 438 1781 497
rect 1707 404 1727 438
rect 1761 404 1781 438
rect 1707 362 1781 404
rect 1707 328 1725 362
rect 1759 328 1781 362
rect 1707 297 1781 328
rect 1811 485 1867 497
rect 1811 451 1822 485
rect 1856 451 1867 485
rect 1811 417 1867 451
rect 1811 383 1822 417
rect 1856 383 1867 417
rect 1811 297 1867 383
rect 1897 436 1950 497
rect 1897 402 1908 436
rect 1942 402 1950 436
rect 1897 362 1950 402
rect 1897 328 1908 362
rect 1942 328 1950 362
rect 1897 297 1950 328
<< ndiffc >>
rect 39 55 73 89
rect 123 107 157 141
rect 208 55 242 89
rect 294 107 328 141
rect 396 55 430 89
rect 482 107 516 141
rect 568 55 602 89
rect 654 107 688 141
rect 752 55 786 89
rect 848 107 882 141
rect 934 55 968 89
rect 1020 107 1054 141
rect 1105 55 1139 89
rect 1217 55 1251 89
rect 1302 123 1336 157
rect 1388 55 1422 89
rect 1474 123 1508 157
rect 1578 85 1612 119
rect 1665 55 1699 89
rect 1751 85 1785 119
rect 1837 55 1871 89
rect 1923 85 1957 119
<< pdiffc >>
rect 36 451 70 485
rect 36 383 70 417
rect 122 379 156 413
rect 122 311 156 345
rect 208 455 242 489
rect 208 387 242 421
rect 294 383 328 417
rect 294 314 328 348
rect 380 455 414 489
rect 380 387 414 421
rect 466 383 500 417
rect 466 315 500 349
rect 552 455 586 489
rect 552 387 586 421
rect 638 383 672 417
rect 638 314 672 348
rect 723 451 757 485
rect 723 383 757 417
rect 829 451 863 485
rect 829 383 863 417
rect 914 383 948 417
rect 914 314 948 348
rect 1000 455 1034 489
rect 1000 387 1034 421
rect 1086 383 1120 417
rect 1086 314 1120 348
rect 1174 439 1208 473
rect 1174 309 1208 343
rect 1260 455 1294 489
rect 1260 361 1294 395
rect 1346 403 1380 437
rect 1346 309 1380 343
rect 1432 455 1466 489
rect 1432 361 1466 395
rect 1532 408 1566 442
rect 1522 309 1556 343
rect 1632 451 1666 485
rect 1632 379 1666 413
rect 1727 404 1761 438
rect 1725 328 1759 362
rect 1822 451 1856 485
rect 1822 383 1856 417
rect 1908 402 1942 436
rect 1908 328 1942 362
<< poly >>
rect 81 249 369 265
rect 81 215 115 249
rect 149 215 183 249
rect 217 215 251 249
rect 285 215 319 249
rect 353 215 369 249
rect 81 199 369 215
rect 411 249 749 265
rect 411 215 427 249
rect 461 215 495 249
rect 529 215 563 249
rect 597 215 631 249
rect 665 215 699 249
rect 733 215 749 249
rect 411 199 749 215
rect 791 249 1161 265
rect 791 215 807 249
rect 841 215 875 249
rect 909 215 943 249
rect 977 215 1011 249
rect 1045 215 1079 249
rect 1113 215 1161 249
rect 791 199 1161 215
rect 1219 249 1549 265
rect 1219 215 1289 249
rect 1323 215 1357 249
rect 1391 215 1425 249
rect 1459 215 1493 249
rect 1527 215 1549 249
rect 1219 199 1549 215
rect 1591 249 1998 265
rect 1591 215 1608 249
rect 1642 215 1676 249
rect 1710 215 1744 249
rect 1778 215 1812 249
rect 1846 215 1880 249
rect 1914 215 1948 249
rect 1982 215 1998 249
rect 1591 199 1998 215
<< polycont >>
rect 115 215 149 249
rect 183 215 217 249
rect 251 215 285 249
rect 319 215 353 249
rect 427 215 461 249
rect 495 215 529 249
rect 563 215 597 249
rect 631 215 665 249
rect 699 215 733 249
rect 807 215 841 249
rect 875 215 909 249
rect 943 215 977 249
rect 1011 215 1045 249
rect 1079 215 1113 249
rect 1289 215 1323 249
rect 1357 215 1391 249
rect 1425 215 1459 249
rect 1493 215 1527 249
rect 1608 215 1642 249
rect 1676 215 1710 249
rect 1744 215 1778 249
rect 1812 215 1846 249
rect 1880 215 1914 249
rect 1948 215 1982 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 1244 489 1310 527
rect 20 485 208 489
rect 20 451 36 485
rect 70 455 208 485
rect 242 455 380 489
rect 414 455 552 489
rect 586 485 774 489
rect 586 455 723 485
rect 70 451 723 455
rect 757 451 774 485
rect 20 417 72 451
rect 206 421 244 451
rect 20 383 36 417
rect 70 383 72 417
rect 20 367 72 383
rect 106 413 172 417
rect 106 379 122 413
rect 156 379 172 413
rect 106 345 172 379
rect 206 387 208 421
rect 242 387 244 421
rect 378 421 416 451
rect 206 371 244 387
rect 278 383 294 417
rect 328 383 344 417
rect 106 331 122 345
rect 29 311 122 331
rect 156 337 172 345
rect 278 348 344 383
rect 378 387 380 421
rect 414 387 416 421
rect 550 421 588 451
rect 378 371 416 387
rect 450 383 466 417
rect 500 383 516 417
rect 278 337 294 348
rect 156 314 294 337
rect 328 314 344 348
rect 156 311 344 314
rect 29 295 344 311
rect 450 349 516 383
rect 550 387 552 421
rect 586 387 588 421
rect 722 417 774 451
rect 550 371 588 387
rect 622 383 638 417
rect 672 383 688 417
rect 450 315 466 349
rect 500 337 516 349
rect 622 348 688 383
rect 722 383 723 417
rect 757 383 774 417
rect 722 367 774 383
rect 812 485 1000 489
rect 812 451 829 485
rect 863 455 1000 485
rect 1034 473 1210 489
rect 1034 455 1174 473
rect 863 451 1036 455
rect 812 417 864 451
rect 998 421 1036 451
rect 812 383 829 417
rect 863 383 864 417
rect 812 367 864 383
rect 898 383 914 417
rect 948 383 964 417
rect 622 337 638 348
rect 500 315 638 337
rect 450 314 638 315
rect 672 331 688 348
rect 898 348 964 383
rect 998 387 1000 421
rect 1034 387 1036 421
rect 1172 439 1174 455
rect 1208 439 1210 473
rect 998 371 1036 387
rect 1070 383 1086 417
rect 1120 383 1136 417
rect 898 331 914 348
rect 672 314 914 331
rect 948 337 964 348
rect 1070 348 1136 383
rect 1070 337 1086 348
rect 948 314 1086 337
rect 1120 314 1136 348
rect 450 295 1136 314
rect 1172 343 1210 439
rect 1244 455 1260 489
rect 1294 455 1310 489
rect 1416 489 1482 527
rect 1244 395 1310 455
rect 1244 361 1260 395
rect 1294 361 1310 395
rect 1244 357 1310 361
rect 1344 437 1382 463
rect 1344 403 1346 437
rect 1380 403 1382 437
rect 1172 309 1174 343
rect 1208 323 1210 343
rect 1344 343 1382 403
rect 1416 455 1432 489
rect 1466 455 1482 489
rect 1616 485 1682 527
rect 1416 395 1482 455
rect 1416 361 1432 395
rect 1466 361 1482 395
rect 1516 442 1582 463
rect 1516 408 1532 442
rect 1566 408 1582 442
rect 1344 323 1346 343
rect 1208 309 1346 323
rect 1380 323 1382 343
rect 1516 343 1582 408
rect 1616 451 1632 485
rect 1666 451 1682 485
rect 1806 485 1872 527
rect 1616 413 1682 451
rect 1616 379 1632 413
rect 1666 379 1682 413
rect 1716 438 1768 458
rect 1716 404 1727 438
rect 1761 404 1768 438
rect 1516 323 1522 343
rect 1380 309 1522 323
rect 1556 333 1582 343
rect 1716 362 1768 404
rect 1806 451 1822 485
rect 1856 451 1872 485
rect 1806 417 1872 451
rect 1806 383 1822 417
rect 1856 383 1872 417
rect 1906 436 1954 452
rect 1906 402 1908 436
rect 1942 402 1954 436
rect 1716 333 1725 362
rect 1556 328 1725 333
rect 1759 334 1768 362
rect 1906 362 1954 402
rect 1906 334 1908 362
rect 1759 328 1908 334
rect 1942 328 1954 362
rect 1556 309 1954 328
rect 29 157 64 295
rect 1172 289 1954 309
rect 99 249 369 255
rect 99 215 115 249
rect 149 215 183 249
rect 217 215 251 249
rect 285 215 319 249
rect 353 215 369 249
rect 99 204 369 215
rect 411 249 749 255
rect 411 215 427 249
rect 461 215 495 249
rect 529 215 563 249
rect 597 215 631 249
rect 665 215 699 249
rect 733 215 749 249
rect 411 204 749 215
rect 791 249 1130 255
rect 791 215 807 249
rect 841 215 875 249
rect 909 215 943 249
rect 977 215 1011 249
rect 1045 215 1079 249
rect 1113 215 1130 249
rect 791 204 1130 215
rect 1219 249 1549 255
rect 1219 215 1289 249
rect 1323 215 1357 249
rect 1391 215 1425 249
rect 1459 215 1493 249
rect 1527 215 1549 249
rect 1219 204 1549 215
rect 1592 249 1998 255
rect 1592 215 1608 249
rect 1642 215 1676 249
rect 1710 215 1744 249
rect 1778 215 1812 249
rect 1846 215 1880 249
rect 1914 215 1948 249
rect 1982 215 1998 249
rect 1592 204 1998 215
rect 29 141 1302 157
rect 29 123 123 141
rect 157 123 294 141
rect 157 107 158 123
rect 123 91 158 107
rect 292 107 294 123
rect 328 123 482 141
rect 328 107 330 123
rect 292 91 330 107
rect 480 107 482 123
rect 516 123 654 141
rect 516 107 518 123
rect 480 91 518 107
rect 652 107 654 123
rect 688 123 848 141
rect 688 107 702 123
rect 652 91 702 107
rect 836 107 848 123
rect 882 123 1020 141
rect 882 107 884 123
rect 836 91 884 107
rect 1018 107 1020 123
rect 1054 123 1302 141
rect 1336 123 1474 157
rect 1508 123 1524 157
rect 1577 123 1973 157
rect 1054 107 1055 123
rect 1018 91 1055 107
rect 1577 119 1615 123
rect 1577 89 1578 119
rect 23 55 39 89
rect 73 55 89 89
rect 23 17 89 55
rect 192 55 208 89
rect 242 55 258 89
rect 192 17 258 55
rect 364 55 396 89
rect 430 55 446 89
rect 364 17 446 55
rect 552 55 568 89
rect 602 55 618 89
rect 552 17 618 55
rect 736 55 752 89
rect 786 55 802 89
rect 736 17 802 55
rect 918 55 934 89
rect 968 55 984 89
rect 918 17 984 55
rect 1089 55 1105 89
rect 1139 55 1156 89
rect 1196 55 1217 89
rect 1251 55 1388 89
rect 1422 85 1578 89
rect 1612 85 1615 119
rect 1749 119 1787 123
rect 1422 55 1615 85
rect 1649 55 1665 89
rect 1699 55 1715 89
rect 1749 85 1751 119
rect 1785 85 1787 119
rect 1921 119 1973 123
rect 1749 60 1787 85
rect 1089 17 1156 55
rect 1649 17 1715 55
rect 1821 55 1837 89
rect 1871 55 1887 89
rect 1921 85 1923 119
rect 1957 85 1973 119
rect 1921 58 1973 85
rect 1821 17 1887 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
<< metal1 >>
rect 0 561 2024 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 0 496 2024 527
rect 0 17 2024 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
rect 0 -48 2024 -17
<< labels >>
flabel locali s 122 221 156 255 0 FreeSans 340 0 0 0 D1
port 5 nsew signal input
flabel locali s 490 221 524 255 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 858 221 892 255 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 1780 221 1814 255 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1228 221 1262 255 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 30 153 64 187 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 a2111oi_4
rlabel metal1 s 0 -48 2024 48 1 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 496 2024 592 1 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2024 544
string GDS_END 3820934
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3806770
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 50.600 0.000 
<< end >>
