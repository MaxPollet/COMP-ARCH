magic
tech sky130A
magscale 1 2
timestamp 1681267127
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 1 21 643 203
rect 30 13 212 21
rect 30 -17 64 13
<< locali >>
rect 18 369 85 485
rect 18 157 72 369
rect 108 193 156 333
rect 192 193 250 333
rect 18 123 258 157
rect 294 151 342 333
rect 378 151 442 333
rect 556 199 617 323
rect 18 57 69 123
rect 224 93 258 123
rect 537 93 603 161
rect 224 59 603 93
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 119 403 169 493
rect 224 439 290 527
rect 352 403 386 493
rect 443 439 509 527
rect 553 403 603 493
rect 119 369 603 403
rect 124 17 190 89
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
rlabel locali s 556 199 617 323 6 A1
port 1 nsew signal input
rlabel locali s 378 151 442 333 6 A2
port 2 nsew signal input
rlabel locali s 294 151 342 333 6 A3
port 3 nsew signal input
rlabel locali s 192 193 250 333 6 A4
port 4 nsew signal input
rlabel locali s 108 193 156 333 6 B1
port 5 nsew signal input
rlabel metal1 s 0 -48 644 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 13 8 VNB
port 7 nsew ground bidirectional
rlabel pwell s 30 13 212 21 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 1 21 643 203 6 VNB
port 7 nsew ground bidirectional
rlabel nwell s -38 261 682 582 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 496 644 592 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 224 59 603 93 6 Y
port 10 nsew signal output
rlabel locali s 537 93 603 161 6 Y
port 10 nsew signal output
rlabel locali s 224 93 258 123 6 Y
port 10 nsew signal output
rlabel locali s 18 57 69 123 6 Y
port 10 nsew signal output
rlabel locali s 18 123 258 157 6 Y
port 10 nsew signal output
rlabel locali s 18 157 72 369 6 Y
port 10 nsew signal output
rlabel locali s 18 369 85 485 6 Y
port 10 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 644 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 3556200
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3549478
<< end >>
