magic
tech sky130A
magscale 1 2
timestamp 1681267127
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 1 67 735 203
rect 1 21 637 67
rect 29 -17 63 21
<< scnmos >>
rect 79 47 109 177
rect 153 47 183 177
rect 267 47 297 177
rect 353 47 383 177
rect 439 47 469 177
rect 525 47 555 177
rect 626 93 656 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 267 297 297 497
rect 357 297 387 497
rect 441 297 471 497
rect 525 297 555 497
rect 626 297 656 381
<< ndiff >>
rect 27 161 79 177
rect 27 127 35 161
rect 69 127 79 161
rect 27 93 79 127
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 47 153 177
rect 183 89 267 177
rect 183 55 207 89
rect 241 55 267 89
rect 183 47 267 55
rect 297 149 353 177
rect 297 115 307 149
rect 341 115 353 149
rect 297 47 353 115
rect 383 89 439 177
rect 383 55 393 89
rect 427 55 439 89
rect 383 47 439 55
rect 469 165 525 177
rect 469 131 480 165
rect 514 131 525 165
rect 469 47 525 131
rect 555 93 626 177
rect 656 153 709 177
rect 656 119 666 153
rect 700 119 709 153
rect 656 93 709 119
rect 555 89 611 93
rect 555 55 565 89
rect 599 55 611 89
rect 555 47 611 55
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 297 79 451
rect 109 349 163 497
rect 109 315 119 349
rect 153 315 163 349
rect 109 297 163 315
rect 193 489 267 497
rect 193 455 214 489
rect 248 455 267 489
rect 193 297 267 455
rect 297 341 357 497
rect 297 307 313 341
rect 347 307 357 341
rect 297 297 357 307
rect 387 489 441 497
rect 387 455 397 489
rect 431 455 441 489
rect 387 297 441 455
rect 471 341 525 497
rect 471 307 481 341
rect 515 307 525 341
rect 471 297 525 307
rect 555 489 611 497
rect 555 455 565 489
rect 599 455 611 489
rect 555 381 611 455
rect 555 297 626 381
rect 656 356 709 381
rect 656 322 667 356
rect 701 322 709 356
rect 656 297 709 322
<< ndiffc >>
rect 35 127 69 161
rect 35 59 69 93
rect 207 55 241 89
rect 307 115 341 149
rect 393 55 427 89
rect 480 131 514 165
rect 666 119 700 153
rect 565 55 599 89
<< pdiffc >>
rect 35 451 69 485
rect 119 315 153 349
rect 214 455 248 489
rect 313 307 347 341
rect 397 455 431 489
rect 481 307 515 341
rect 565 455 599 489
rect 667 322 701 356
<< poly >>
rect 33 249 109 265
rect 33 215 51 249
rect 85 215 109 249
rect 33 199 109 215
rect 151 249 205 265
rect 151 215 161 249
rect 195 215 205 249
rect 151 199 205 215
rect 267 249 555 265
rect 267 215 282 249
rect 316 215 350 249
rect 384 215 418 249
rect 452 215 555 249
rect 267 199 555 215
rect 597 249 656 268
rect 597 215 607 249
rect 641 215 656 249
rect 597 199 656 215
<< polycont >>
rect 51 215 85 249
rect 161 215 195 249
rect 282 215 316 249
rect 350 215 384 249
rect 418 215 452 249
rect 607 215 641 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 18 485 85 527
rect 18 451 35 485
rect 69 451 85 485
rect 198 489 264 527
rect 198 455 214 489
rect 248 455 264 489
rect 381 489 447 527
rect 381 455 397 489
rect 431 455 447 489
rect 549 489 615 527
rect 549 455 565 489
rect 599 455 615 489
rect 33 383 701 417
rect 33 265 67 383
rect 667 356 701 383
rect 103 315 119 349
rect 153 315 263 349
rect 103 300 263 315
rect 297 341 546 349
rect 297 307 313 341
rect 347 307 481 341
rect 515 307 546 341
rect 222 297 263 300
rect 222 287 264 297
rect 229 271 264 287
rect 33 249 85 265
rect 33 215 51 249
rect 33 199 85 215
rect 122 249 195 265
rect 122 215 161 249
rect 122 199 195 215
rect 229 249 452 271
rect 229 215 282 249
rect 316 215 350 249
rect 384 215 418 249
rect 229 199 452 215
rect 229 161 271 199
rect 488 165 546 307
rect 18 127 35 161
rect 69 127 271 161
rect 18 123 271 127
rect 305 149 480 165
rect 18 93 85 123
rect 305 115 307 149
rect 341 131 480 149
rect 514 131 546 165
rect 341 123 546 131
rect 580 265 631 349
rect 701 322 709 340
rect 667 306 709 322
rect 580 249 641 265
rect 580 215 607 249
rect 580 199 641 215
rect 580 125 631 199
rect 675 169 709 306
rect 666 153 709 169
rect 341 115 343 123
rect 305 99 343 115
rect 700 135 709 153
rect 666 99 700 119
rect 18 59 35 93
rect 69 59 85 93
rect 18 51 85 59
rect 191 55 207 89
rect 241 55 257 89
rect 191 17 257 55
rect 377 55 393 89
rect 427 55 443 89
rect 377 17 443 55
rect 549 55 565 89
rect 599 55 615 89
rect 549 17 615 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
flabel locali s 122 221 156 255 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 488 153 522 187 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 580 221 614 255 0 FreeSans 400 0 0 0 A_N
port 1 nsew signal input
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 and2b_4
rlabel metal1 s 0 -48 736 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 736 592 1 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 736 544
string GDS_END 3871442
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3865784
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 18.400 0.000 
<< end >>
