magic
tech sky130A
magscale 1 2
timestamp 1681267127
<< nwell >>
rect -38 261 2430 582
<< pwell >>
rect 1924 201 2391 203
rect 782 157 1236 201
rect 1557 157 2391 201
rect 1 21 2391 157
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 131
rect 163 47 193 131
rect 351 47 381 131
rect 446 47 476 119
rect 552 47 582 119
rect 648 47 678 131
rect 758 47 788 131
rect 858 47 888 175
rect 942 47 972 175
rect 1130 47 1160 175
rect 1225 47 1255 119
rect 1334 47 1364 119
rect 1429 47 1459 131
rect 1515 47 1545 131
rect 1633 47 1663 175
rect 1717 47 1747 175
rect 1905 47 1935 131
rect 2000 47 2030 177
rect 2188 47 2218 131
rect 2283 47 2313 177
<< scpmoshvt >>
rect 79 363 109 491
rect 163 363 193 491
rect 351 413 381 497
rect 444 413 474 497
rect 528 413 558 497
rect 648 413 678 497
rect 754 413 784 497
rect 862 329 892 497
rect 946 329 976 497
rect 1083 329 1113 497
rect 1227 413 1257 497
rect 1311 413 1341 497
rect 1429 413 1459 497
rect 1537 413 1567 497
rect 1633 329 1663 497
rect 1705 329 1735 497
rect 1903 301 1933 429
rect 2000 297 2030 497
rect 2188 353 2218 481
rect 2283 297 2313 497
<< ndiff >>
rect 808 131 858 175
rect 27 119 79 131
rect 27 85 35 119
rect 69 85 79 119
rect 27 47 79 85
rect 109 93 163 131
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 119 245 131
rect 193 85 203 119
rect 237 85 245 119
rect 193 47 245 85
rect 299 93 351 131
rect 299 59 307 93
rect 341 59 351 93
rect 299 47 351 59
rect 381 119 431 131
rect 597 119 648 131
rect 381 111 446 119
rect 381 77 391 111
rect 425 77 446 111
rect 381 47 446 77
rect 476 93 552 119
rect 476 59 497 93
rect 531 59 552 93
rect 476 47 552 59
rect 582 47 648 119
rect 678 89 758 131
rect 678 55 714 89
rect 748 55 758 89
rect 678 47 758 55
rect 788 109 858 131
rect 788 75 798 109
rect 832 75 858 109
rect 788 47 858 75
rect 888 153 942 175
rect 888 119 898 153
rect 932 119 942 153
rect 888 47 942 119
rect 972 127 1024 175
rect 972 93 982 127
rect 1016 93 1024 127
rect 972 47 1024 93
rect 1078 93 1130 175
rect 1078 59 1086 93
rect 1120 59 1130 93
rect 1078 47 1130 59
rect 1160 119 1210 175
rect 1583 131 1633 175
rect 1379 119 1429 131
rect 1160 47 1225 119
rect 1255 93 1334 119
rect 1255 59 1280 93
rect 1314 59 1334 93
rect 1255 47 1334 59
rect 1364 47 1429 119
rect 1459 89 1515 131
rect 1459 55 1471 89
rect 1505 55 1515 89
rect 1459 47 1515 55
rect 1545 109 1633 131
rect 1545 75 1573 109
rect 1607 75 1633 109
rect 1545 47 1633 75
rect 1663 153 1717 175
rect 1663 119 1673 153
rect 1707 119 1717 153
rect 1663 47 1717 119
rect 1747 101 1799 175
rect 1950 131 2000 177
rect 1747 67 1757 101
rect 1791 67 1799 101
rect 1747 47 1799 67
rect 1853 103 1905 131
rect 1853 69 1861 103
rect 1895 69 1905 103
rect 1853 47 1905 69
rect 1935 93 2000 131
rect 1935 59 1956 93
rect 1990 59 2000 93
rect 1935 47 2000 59
rect 2030 127 2082 177
rect 2233 131 2283 177
rect 2030 93 2040 127
rect 2074 93 2082 127
rect 2030 47 2082 93
rect 2136 119 2188 131
rect 2136 85 2144 119
rect 2178 85 2188 119
rect 2136 47 2188 85
rect 2218 93 2283 131
rect 2218 59 2239 93
rect 2273 59 2283 93
rect 2218 47 2283 59
rect 2313 129 2365 177
rect 2313 95 2323 129
rect 2357 95 2365 129
rect 2313 47 2365 95
<< pdiff >>
rect 27 477 79 491
rect 27 443 35 477
rect 69 443 79 477
rect 27 409 79 443
rect 27 375 35 409
rect 69 375 79 409
rect 27 363 79 375
rect 109 461 163 491
rect 109 427 119 461
rect 153 427 163 461
rect 109 363 163 427
rect 193 477 245 491
rect 193 443 203 477
rect 237 443 245 477
rect 193 409 245 443
rect 299 461 351 497
rect 299 427 307 461
rect 341 427 351 461
rect 299 413 351 427
rect 381 477 444 497
rect 381 443 391 477
rect 425 443 444 477
rect 381 413 444 443
rect 474 484 528 497
rect 474 450 484 484
rect 518 450 528 484
rect 474 413 528 450
rect 558 413 648 497
rect 678 475 754 497
rect 678 441 698 475
rect 732 441 754 475
rect 678 413 754 441
rect 784 459 862 497
rect 784 425 818 459
rect 852 425 862 459
rect 784 413 862 425
rect 193 375 203 409
rect 237 375 245 409
rect 800 391 862 413
rect 193 363 245 375
rect 800 357 818 391
rect 852 357 862 391
rect 800 329 862 357
rect 892 329 946 497
rect 976 485 1083 497
rect 976 451 992 485
rect 1026 451 1083 485
rect 976 417 1083 451
rect 976 383 992 417
rect 1026 383 1083 417
rect 976 329 1083 383
rect 1113 413 1227 497
rect 1257 484 1311 497
rect 1257 450 1267 484
rect 1301 450 1311 484
rect 1257 413 1311 450
rect 1341 413 1429 497
rect 1459 485 1537 497
rect 1459 451 1481 485
rect 1515 451 1537 485
rect 1459 413 1537 451
rect 1567 459 1633 497
rect 1567 425 1589 459
rect 1623 425 1633 459
rect 1567 413 1633 425
rect 1113 329 1165 413
rect 1582 329 1633 413
rect 1663 329 1705 497
rect 1735 485 1787 497
rect 1735 451 1745 485
rect 1779 451 1787 485
rect 1735 329 1787 451
rect 1948 485 2000 497
rect 1948 451 1956 485
rect 1990 451 2000 485
rect 1948 429 2000 451
rect 1851 349 1903 429
rect 1851 315 1859 349
rect 1893 315 1903 349
rect 1851 301 1903 315
rect 1933 301 2000 429
rect 1950 297 2000 301
rect 2030 448 2082 497
rect 2233 481 2283 497
rect 2030 414 2040 448
rect 2074 414 2082 448
rect 2030 380 2082 414
rect 2030 346 2040 380
rect 2074 346 2082 380
rect 2136 467 2188 481
rect 2136 433 2144 467
rect 2178 433 2188 467
rect 2136 399 2188 433
rect 2136 365 2144 399
rect 2178 365 2188 399
rect 2136 353 2188 365
rect 2218 473 2283 481
rect 2218 439 2239 473
rect 2273 439 2283 473
rect 2218 405 2283 439
rect 2218 371 2239 405
rect 2273 371 2283 405
rect 2218 353 2283 371
rect 2030 297 2082 346
rect 2233 297 2283 353
rect 2313 449 2365 497
rect 2313 415 2323 449
rect 2357 415 2365 449
rect 2313 381 2365 415
rect 2313 347 2323 381
rect 2357 347 2365 381
rect 2313 297 2365 347
<< ndiffc >>
rect 35 85 69 119
rect 119 59 153 93
rect 203 85 237 119
rect 307 59 341 93
rect 391 77 425 111
rect 497 59 531 93
rect 714 55 748 89
rect 798 75 832 109
rect 898 119 932 153
rect 982 93 1016 127
rect 1086 59 1120 93
rect 1280 59 1314 93
rect 1471 55 1505 89
rect 1573 75 1607 109
rect 1673 119 1707 153
rect 1757 67 1791 101
rect 1861 69 1895 103
rect 1956 59 1990 93
rect 2040 93 2074 127
rect 2144 85 2178 119
rect 2239 59 2273 93
rect 2323 95 2357 129
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 119 427 153 461
rect 203 443 237 477
rect 307 427 341 461
rect 391 443 425 477
rect 484 450 518 484
rect 698 441 732 475
rect 818 425 852 459
rect 203 375 237 409
rect 818 357 852 391
rect 992 451 1026 485
rect 992 383 1026 417
rect 1267 450 1301 484
rect 1481 451 1515 485
rect 1589 425 1623 459
rect 1745 451 1779 485
rect 1956 451 1990 485
rect 1859 315 1893 349
rect 2040 414 2074 448
rect 2040 346 2074 380
rect 2144 433 2178 467
rect 2144 365 2178 399
rect 2239 439 2273 473
rect 2239 371 2273 405
rect 2323 415 2357 449
rect 2323 347 2357 381
<< poly >>
rect 516 365 582 375
rect 516 331 532 365
rect 566 331 582 365
rect 516 321 582 331
rect 648 365 712 381
rect 648 331 668 365
rect 702 331 712 365
rect 648 315 712 331
rect 1203 365 1257 381
rect 1203 331 1213 365
rect 1247 331 1257 365
rect 1203 315 1257 331
rect 1299 365 1365 375
rect 1299 331 1315 365
rect 1349 331 1365 365
rect 1299 321 1365 331
rect 1429 365 1495 381
rect 1429 331 1451 365
rect 1485 331 1495 365
rect 1429 315 1495 331
rect 826 281 892 297
rect 21 264 76 280
rect 21 230 32 264
rect 66 230 76 264
rect 21 214 76 230
rect 118 264 193 274
rect 118 230 134 264
rect 168 230 193 264
rect 118 220 193 230
rect 340 251 394 267
rect 340 217 350 251
rect 384 217 394 251
rect 826 247 836 281
rect 870 247 892 281
rect 826 231 892 247
rect 942 281 1032 297
rect 1717 281 1801 297
rect 942 247 988 281
rect 1022 247 1032 281
rect 1609 265 1663 281
rect 942 231 1032 247
rect 1106 247 1160 263
rect 340 201 394 217
rect 446 191 510 207
rect 446 157 466 191
rect 500 157 510 191
rect 446 141 510 157
rect 552 203 606 219
rect 552 169 562 203
rect 596 169 606 203
rect 552 153 606 169
rect 724 213 784 229
rect 724 179 734 213
rect 768 179 784 213
rect 1106 213 1116 247
rect 1150 213 1160 247
rect 1609 231 1619 265
rect 1653 231 1663 265
rect 1717 247 1757 281
rect 1791 247 1801 281
rect 1717 231 1801 247
rect 1872 253 1936 269
rect 1106 197 1160 213
rect 1501 213 1567 229
rect 1609 215 1663 231
rect 1872 219 1888 253
rect 1922 219 1936 253
rect 724 163 784 179
rect 1225 191 1292 207
rect 1225 157 1248 191
rect 1282 157 1292 191
rect 1501 179 1511 213
rect 1545 179 1567 213
rect 1872 203 1936 219
rect 1978 249 2192 259
rect 1978 215 1988 249
rect 2022 215 2192 249
rect 1978 205 2192 215
rect 2254 249 2313 265
rect 2254 215 2264 249
rect 2298 215 2313 249
rect 2254 199 2313 215
rect 1501 163 1567 179
rect 1225 141 1292 157
<< polycont >>
rect 532 331 566 365
rect 668 331 702 365
rect 1213 331 1247 365
rect 1315 331 1349 365
rect 1451 331 1485 365
rect 32 230 66 264
rect 134 230 168 264
rect 350 217 384 251
rect 836 247 870 281
rect 988 247 1022 281
rect 466 157 500 191
rect 562 169 596 203
rect 734 179 768 213
rect 1116 213 1150 247
rect 1619 231 1653 265
rect 1757 247 1791 281
rect 1888 219 1922 253
rect 1248 157 1282 191
rect 1511 179 1545 213
rect 1988 215 2022 249
rect 2264 215 2298 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2392 561
rect 17 477 69 493
rect 17 443 35 477
rect 17 409 69 443
rect 103 461 169 527
rect 103 427 119 461
rect 153 427 169 461
rect 203 477 248 493
rect 237 443 248 477
rect 17 375 35 409
rect 203 409 248 443
rect 287 461 357 527
rect 287 427 307 461
rect 341 427 357 461
rect 391 477 425 493
rect 468 450 484 484
rect 518 450 634 484
rect 69 391 168 393
rect 69 375 122 391
rect 17 359 122 375
rect 156 357 168 391
rect 17 264 88 325
rect 17 230 32 264
rect 66 230 88 264
rect 17 195 88 230
rect 122 264 168 357
rect 122 230 134 264
rect 122 161 168 230
rect 17 127 168 161
rect 237 375 248 409
rect 391 393 425 443
rect 203 187 248 375
rect 203 153 214 187
rect 17 119 69 127
rect 17 85 35 119
rect 203 119 248 153
rect 282 359 425 393
rect 282 165 316 359
rect 466 357 490 391
rect 524 365 566 391
rect 524 357 532 365
rect 466 331 532 357
rect 350 251 432 325
rect 384 217 432 251
rect 350 201 432 217
rect 466 315 566 331
rect 466 191 510 315
rect 600 281 634 450
rect 682 475 758 527
rect 976 485 1042 527
rect 682 441 698 475
rect 732 441 758 475
rect 818 459 852 475
rect 818 407 852 425
rect 976 451 992 485
rect 1026 451 1042 485
rect 1465 485 1541 527
rect 976 417 1042 451
rect 1251 450 1267 484
rect 1301 450 1417 484
rect 1465 451 1481 485
rect 1515 451 1541 485
rect 1729 485 2006 527
rect 1589 459 1623 475
rect 668 391 938 407
rect 668 365 818 391
rect 702 357 818 365
rect 852 357 938 391
rect 976 383 992 417
rect 1026 383 1042 417
rect 1213 391 1260 397
rect 702 331 718 357
rect 668 315 718 331
rect 820 281 870 297
rect 600 247 836 281
rect 600 239 680 247
rect 282 127 425 165
rect 500 157 510 191
rect 466 141 510 157
rect 546 169 562 203
rect 596 187 612 203
rect 546 153 578 169
rect 546 129 612 153
rect 17 69 69 85
rect 103 59 119 93
rect 153 59 169 93
rect 237 85 248 119
rect 391 111 425 127
rect 203 69 248 85
rect 103 17 169 59
rect 287 59 307 93
rect 341 59 357 93
rect 646 93 680 239
rect 826 231 870 247
rect 904 213 938 357
rect 1213 365 1226 391
rect 1247 331 1260 357
rect 972 323 1173 331
rect 972 289 1134 323
rect 1168 289 1173 323
rect 1213 315 1260 331
rect 1308 365 1349 381
rect 1308 331 1315 365
rect 972 283 1173 289
rect 972 281 1038 283
rect 972 247 988 281
rect 1022 247 1038 281
rect 1308 261 1349 331
rect 1225 255 1349 261
rect 1100 213 1116 247
rect 1150 213 1166 247
rect 718 179 734 213
rect 768 193 784 213
rect 768 187 800 193
rect 718 153 766 179
rect 904 179 1166 213
rect 1225 221 1226 255
rect 1260 225 1349 255
rect 1383 281 1417 450
rect 1729 451 1745 485
rect 1779 451 1956 485
rect 1990 451 2006 485
rect 1589 417 1623 425
rect 2040 448 2097 493
rect 1451 383 2006 417
rect 1451 365 1501 383
rect 1485 331 1501 365
rect 1451 315 1501 331
rect 1383 265 1653 281
rect 1383 247 1619 265
rect 1260 221 1282 225
rect 1225 191 1282 221
rect 904 153 948 179
rect 718 147 800 153
rect 882 119 898 153
rect 932 119 948 153
rect 1225 157 1248 191
rect 982 127 1016 143
rect 1225 141 1282 157
rect 391 61 425 77
rect 287 17 357 59
rect 481 59 497 93
rect 531 59 680 93
rect 481 53 680 59
rect 714 89 748 105
rect 714 17 748 55
rect 782 75 798 109
rect 832 85 848 109
rect 1383 93 1417 247
rect 1609 231 1619 247
rect 1609 215 1653 231
rect 1492 187 1511 213
rect 1492 153 1502 187
rect 1545 179 1567 213
rect 1536 153 1567 179
rect 1687 156 1723 383
rect 1492 147 1567 153
rect 1657 153 1723 156
rect 1657 119 1673 153
rect 1707 119 1723 153
rect 1757 323 1859 349
rect 1757 289 1778 323
rect 1812 315 1859 323
rect 1893 315 1909 349
rect 1757 281 1812 289
rect 1791 247 1812 281
rect 1972 265 2006 383
rect 2074 414 2097 448
rect 2040 380 2097 414
rect 2074 346 2097 380
rect 2040 326 2097 346
rect 1757 185 1812 247
rect 1863 253 1938 265
rect 1863 219 1888 253
rect 1922 219 1938 253
rect 1972 249 2022 265
rect 1972 215 1988 249
rect 1972 199 2022 215
rect 1757 151 1895 185
rect 982 85 1016 93
rect 832 75 1016 85
rect 782 51 1016 75
rect 1070 59 1086 93
rect 1120 59 1136 93
rect 1070 17 1136 59
rect 1264 59 1280 93
rect 1314 59 1417 93
rect 1264 53 1417 59
rect 1453 89 1505 105
rect 1453 55 1471 89
rect 1453 17 1505 55
rect 1557 75 1573 109
rect 1607 85 1623 109
rect 1757 101 1791 117
rect 1607 75 1757 85
rect 1557 67 1757 75
rect 1557 51 1791 67
rect 1848 103 1895 151
rect 1848 69 1861 103
rect 1848 53 1895 69
rect 1940 93 2006 161
rect 2056 143 2097 326
rect 1940 59 1956 93
rect 1990 59 2006 93
rect 1940 17 2006 59
rect 2040 127 2097 143
rect 2074 93 2097 127
rect 2040 51 2097 93
rect 2131 467 2194 483
rect 2131 433 2144 467
rect 2178 433 2194 467
rect 2131 399 2194 433
rect 2131 365 2144 399
rect 2178 365 2194 399
rect 2131 265 2194 365
rect 2230 473 2289 527
rect 2230 439 2239 473
rect 2273 439 2289 473
rect 2230 405 2289 439
rect 2230 371 2239 405
rect 2273 371 2289 405
rect 2230 353 2289 371
rect 2323 449 2375 493
rect 2357 415 2375 449
rect 2323 381 2375 415
rect 2357 347 2375 381
rect 2323 289 2375 347
rect 2131 249 2298 265
rect 2131 215 2264 249
rect 2131 199 2298 215
rect 2131 119 2194 199
rect 2332 165 2375 289
rect 2131 85 2144 119
rect 2178 85 2194 119
rect 2323 129 2375 165
rect 2131 51 2194 85
rect 2230 93 2289 109
rect 2230 59 2239 93
rect 2273 59 2289 93
rect 2230 17 2289 59
rect 2357 95 2375 129
rect 2323 51 2375 95
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2392 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 122 357 156 391
rect 214 153 248 187
rect 490 357 524 391
rect 578 169 596 187
rect 596 169 612 187
rect 578 153 612 169
rect 1226 365 1260 391
rect 1226 357 1247 365
rect 1247 357 1260 365
rect 1134 289 1168 323
rect 766 179 768 187
rect 768 179 800 187
rect 766 153 800 179
rect 1226 221 1260 255
rect 1502 179 1511 187
rect 1511 179 1536 187
rect 1502 153 1536 179
rect 1778 289 1812 323
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
<< metal1 >>
rect 0 561 2392 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2392 561
rect 0 496 2392 527
rect 110 391 168 397
rect 110 357 122 391
rect 156 388 168 391
rect 478 391 536 397
rect 478 388 490 391
rect 156 360 490 388
rect 156 357 168 360
rect 110 351 168 357
rect 478 357 490 360
rect 524 388 536 391
rect 1214 391 1272 397
rect 1214 388 1226 391
rect 524 360 1226 388
rect 524 357 536 360
rect 478 351 536 357
rect 1214 357 1226 360
rect 1260 357 1272 391
rect 1214 351 1272 357
rect 1122 323 1180 329
rect 1122 289 1134 323
rect 1168 320 1180 323
rect 1766 323 1824 329
rect 1766 320 1778 323
rect 1168 292 1778 320
rect 1168 289 1180 292
rect 1122 283 1180 289
rect 1766 289 1778 292
rect 1812 289 1824 323
rect 1766 283 1824 289
rect 1214 255 1272 261
rect 1214 252 1226 255
rect 585 224 1226 252
rect 585 193 624 224
rect 1214 221 1226 224
rect 1260 221 1272 255
rect 1214 215 1272 221
rect 202 187 260 193
rect 202 153 214 187
rect 248 184 260 187
rect 566 187 624 193
rect 566 184 578 187
rect 248 156 578 184
rect 248 153 260 156
rect 202 147 260 153
rect 566 153 578 156
rect 612 153 624 187
rect 566 147 624 153
rect 754 187 812 193
rect 754 153 766 187
rect 800 184 812 187
rect 1490 187 1548 193
rect 1490 184 1502 187
rect 800 156 1502 184
rect 800 153 812 156
rect 754 147 812 153
rect 1490 153 1502 156
rect 1536 153 1548 187
rect 1490 147 1548 153
rect 0 17 2392 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2392 17
rect 0 -48 2392 -17
<< labels >>
flabel locali s 1863 219 1938 265 0 FreeSans 400 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 30 -17 64 17 3 FreeSans 400 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel locali s 30 221 64 255 0 FreeSans 400 0 0 0 CLK
port 1 nsew clock input
flabel locali s 30 289 64 323 0 FreeSans 400 0 0 0 CLK
port 1 nsew clock input
flabel locali s 766 153 800 187 0 FreeSans 400 0 0 0 SET_B
port 4 nsew signal input
flabel locali s 2328 85 2362 119 0 FreeSans 400 0 0 0 Q
port 9 nsew signal output
flabel locali s 2328 357 2362 391 0 FreeSans 400 0 0 0 Q
port 9 nsew signal output
flabel locali s 2328 425 2362 459 0 FreeSans 400 0 0 0 Q
port 9 nsew signal output
flabel locali s 30 527 64 561 3 FreeSans 400 0 0 0 VPWR
port 8 nsew power bidirectional abutment
flabel locali s 398 221 432 255 0 FreeSans 200 0 0 0 D
port 2 nsew signal input
flabel locali s 398 289 432 323 0 FreeSans 200 0 0 0 D
port 2 nsew signal input
flabel locali s 2048 425 2082 459 0 FreeSans 400 0 0 0 Q_N
port 10 nsew signal output
flabel locali s 2048 357 2082 391 0 FreeSans 400 0 0 0 Q_N
port 10 nsew signal output
flabel locali s 2048 85 2082 119 0 FreeSans 400 0 0 0 Q_N
port 10 nsew signal output
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
flabel nwell s 30 527 64 561 3 FreeSans 400 0 0 0 VPB
port 7 nsew power bidirectional
flabel nwell s 47 544 47 544 0 FreeSans 200 0 0 0 VPB
flabel pwell s 30 -17 64 17 3 FreeSans 400 0 0 0 VNB
port 6 nsew ground bidirectional
flabel pwell s 47 0 47 0 0 FreeSans 200 0 0 0 VNB
rlabel comment s 0 0 0 0 4 dfbbp_1
rlabel locali s 1492 147 1567 213 1 SET_B
port 4 nsew signal input
rlabel metal1 s 1490 184 1548 193 1 SET_B
port 4 nsew signal input
rlabel metal1 s 1490 147 1548 156 1 SET_B
port 4 nsew signal input
rlabel metal1 s 754 184 812 193 1 SET_B
port 4 nsew signal input
rlabel metal1 s 754 156 1548 184 1 SET_B
port 4 nsew signal input
rlabel metal1 s 754 147 812 156 1 SET_B
port 4 nsew signal input
rlabel metal1 s 0 -48 2392 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 2392 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2392 544
string GDS_END 3423836
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3404818
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
