magic
tech sky130A
magscale 1 2
timestamp 1681267127
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 1 163 187 203
rect 453 163 643 203
rect 1 67 643 163
rect 30 27 643 67
rect 30 -17 64 27
rect 456 21 643 27
<< scnmos >>
rect 79 93 109 177
rect 266 53 296 137
rect 338 53 368 137
rect 419 53 449 137
rect 535 47 565 177
<< scpmoshvt >>
rect 79 413 109 497
rect 261 311 291 395
rect 345 311 375 395
rect 440 297 470 381
rect 535 297 565 497
<< ndiff >>
rect 27 163 79 177
rect 27 129 35 163
rect 69 129 79 163
rect 27 93 79 129
rect 109 165 161 177
rect 109 131 119 165
rect 153 131 161 165
rect 479 137 535 177
rect 109 120 161 131
rect 109 93 159 120
rect 216 110 266 137
rect 215 109 266 110
rect 214 99 266 109
rect 214 65 222 99
rect 256 65 266 99
rect 214 53 266 65
rect 296 53 338 137
rect 368 53 419 137
rect 449 109 535 137
rect 449 75 491 109
rect 525 75 535 109
rect 449 53 535 75
rect 482 47 535 53
rect 565 119 617 177
rect 565 85 575 119
rect 609 85 617 119
rect 565 47 617 85
<< pdiff >>
rect 27 475 79 497
rect 27 441 35 475
rect 69 441 79 475
rect 27 413 79 441
rect 109 469 161 497
rect 109 435 119 469
rect 153 435 161 469
rect 109 423 161 435
rect 483 485 535 497
rect 483 451 491 485
rect 525 451 535 485
rect 483 438 535 451
rect 109 413 159 423
rect 211 381 261 395
rect 209 369 261 381
rect 209 335 217 369
rect 251 335 261 369
rect 209 311 261 335
rect 291 387 345 395
rect 291 353 301 387
rect 335 353 345 387
rect 291 311 345 353
rect 375 381 425 395
rect 485 381 535 438
rect 375 362 440 381
rect 375 328 395 362
rect 429 328 440 362
rect 375 311 440 328
rect 390 297 440 311
rect 470 297 535 381
rect 565 471 617 497
rect 565 437 575 471
rect 609 437 617 471
rect 565 403 617 437
rect 565 369 575 403
rect 609 369 617 403
rect 565 297 617 369
<< ndiffc >>
rect 35 129 69 163
rect 119 131 153 165
rect 222 65 256 99
rect 491 75 525 109
rect 575 85 609 119
<< pdiffc >>
rect 35 441 69 475
rect 119 435 153 469
rect 491 451 525 485
rect 217 335 251 369
rect 301 353 335 387
rect 395 328 429 362
rect 575 437 609 471
rect 575 369 609 403
<< poly >>
rect 345 477 402 500
rect 345 443 358 477
rect 392 443 402 477
rect 345 427 402 443
rect 22 323 109 339
rect 22 289 35 323
rect 69 289 109 323
rect 22 249 109 289
rect 22 215 35 249
rect 69 215 109 249
rect 22 199 109 215
rect 212 249 296 265
rect 212 215 222 249
rect 256 215 296 249
rect 212 199 296 215
rect 419 249 473 265
rect 419 215 429 249
rect 463 215 473 249
rect 419 199 473 215
rect 515 249 569 265
rect 515 215 525 249
rect 559 215 569 249
rect 515 199 569 215
<< polycont >>
rect 358 443 392 477
rect 35 289 69 323
rect 35 215 69 249
rect 222 215 256 249
rect 429 215 463 249
rect 525 215 559 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 17 475 69 527
rect 17 441 35 475
rect 17 425 69 441
rect 119 469 153 493
rect 17 323 85 391
rect 17 289 35 323
rect 69 289 85 323
rect 17 249 85 289
rect 17 215 35 249
rect 69 215 85 249
rect 119 249 153 435
rect 201 426 324 527
rect 201 369 251 392
rect 201 335 217 369
rect 285 391 324 426
rect 358 477 453 493
rect 392 443 453 477
rect 358 425 453 443
rect 487 485 530 527
rect 487 451 491 485
rect 525 451 530 485
rect 487 418 530 451
rect 572 471 627 493
rect 572 437 575 471
rect 609 437 627 471
rect 572 403 627 437
rect 285 387 351 391
rect 285 353 301 387
rect 335 353 351 387
rect 395 362 538 378
rect 201 319 251 335
rect 429 328 538 362
rect 572 369 575 403
rect 609 369 627 403
rect 572 353 627 369
rect 395 319 538 328
rect 201 285 559 319
rect 119 215 222 249
rect 256 215 278 249
rect 119 199 278 215
rect 119 181 169 199
rect 17 163 69 181
rect 17 129 35 163
rect 17 17 69 129
rect 103 165 169 181
rect 103 131 119 165
rect 153 131 169 165
rect 103 97 169 131
rect 312 114 363 285
rect 513 249 559 285
rect 205 99 363 114
rect 205 65 222 99
rect 256 65 363 99
rect 205 61 363 65
rect 397 215 429 249
rect 463 215 479 249
rect 397 145 479 215
rect 513 215 525 249
rect 513 199 559 215
rect 593 147 627 353
rect 397 61 437 145
rect 575 119 627 147
rect 475 75 491 109
rect 525 75 541 109
rect 475 17 541 75
rect 609 85 627 119
rect 575 51 627 85
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
flabel locali s 30 289 64 323 0 FreeSans 400 0 0 0 A_N
port 1 nsew signal input
flabel locali s 397 425 431 459 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel locali s 581 425 615 459 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel locali s 397 153 431 187 0 FreeSans 400 0 0 0 C
port 3 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 400 0 0 0 A_N
port 1 nsew signal input
flabel locali s 580 85 614 119 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel locali s 30 357 64 391 0 FreeSans 400 0 0 0 A_N
port 1 nsew signal input
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 and3b_1
rlabel metal1 s 0 -48 644 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 644 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 644 544
string GDS_END 3877840
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3871498
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 16.100 0.000 
<< end >>
