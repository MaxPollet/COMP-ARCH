magic
tech sky130A
magscale 1 2
timestamp 1681267127
<< nwell >>
rect -38 261 1142 582
<< pwell >>
rect 825 157 1103 203
rect 1 21 1103 157
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 131
rect 163 47 193 131
rect 351 47 381 131
rect 435 47 465 131
rect 530 47 560 119
rect 620 47 650 119
rect 715 47 745 131
rect 903 47 933 177
rect 995 47 1025 177
<< scpmoshvt >>
rect 79 363 109 491
rect 163 363 193 491
rect 351 369 381 497
rect 435 369 465 497
rect 530 413 560 497
rect 614 413 644 497
rect 715 413 745 497
rect 903 297 933 497
rect 995 297 1025 497
<< ndiff >>
rect 27 119 79 131
rect 27 85 35 119
rect 69 85 79 119
rect 27 47 79 85
rect 109 93 163 131
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 119 245 131
rect 193 85 203 119
rect 237 85 245 119
rect 193 47 245 85
rect 299 119 351 131
rect 299 85 307 119
rect 341 85 351 119
rect 299 47 351 85
rect 381 89 435 131
rect 381 55 391 89
rect 425 55 435 89
rect 381 47 435 55
rect 465 119 515 131
rect 665 119 715 131
rect 465 47 530 119
rect 560 107 620 119
rect 560 73 570 107
rect 604 73 620 107
rect 560 47 620 73
rect 650 47 715 119
rect 745 93 797 131
rect 745 59 755 93
rect 789 59 797 93
rect 745 47 797 59
rect 851 102 903 177
rect 851 68 859 102
rect 893 68 903 102
rect 851 47 903 68
rect 933 127 995 177
rect 933 93 951 127
rect 985 93 995 127
rect 933 47 995 93
rect 1025 133 1077 177
rect 1025 99 1035 133
rect 1069 99 1077 133
rect 1025 47 1077 99
<< pdiff >>
rect 27 477 79 491
rect 27 443 35 477
rect 69 443 79 477
rect 27 409 79 443
rect 27 375 35 409
rect 69 375 79 409
rect 27 363 79 375
rect 109 461 163 491
rect 109 427 119 461
rect 153 427 163 461
rect 109 363 163 427
rect 193 477 245 491
rect 193 443 203 477
rect 237 443 245 477
rect 193 409 245 443
rect 193 375 203 409
rect 237 375 245 409
rect 193 363 245 375
rect 299 483 351 497
rect 299 449 307 483
rect 341 449 351 483
rect 299 415 351 449
rect 299 381 307 415
rect 341 381 351 415
rect 299 369 351 381
rect 381 485 435 497
rect 381 451 391 485
rect 425 451 435 485
rect 381 417 435 451
rect 381 383 391 417
rect 425 383 435 417
rect 381 369 435 383
rect 465 413 530 497
rect 560 485 614 497
rect 560 451 570 485
rect 604 451 614 485
rect 560 413 614 451
rect 644 413 715 497
rect 745 485 797 497
rect 745 451 755 485
rect 789 451 797 485
rect 745 413 797 451
rect 851 471 903 497
rect 851 437 859 471
rect 893 437 903 471
rect 465 369 515 413
rect 851 368 903 437
rect 851 334 859 368
rect 893 334 903 368
rect 851 297 903 334
rect 933 484 995 497
rect 933 450 951 484
rect 985 450 995 484
rect 933 364 995 450
rect 933 330 951 364
rect 985 330 995 364
rect 933 297 995 330
rect 1025 475 1077 497
rect 1025 441 1035 475
rect 1069 441 1077 475
rect 1025 384 1077 441
rect 1025 350 1035 384
rect 1069 350 1077 384
rect 1025 297 1077 350
<< ndiffc >>
rect 35 85 69 119
rect 119 59 153 93
rect 203 85 237 119
rect 307 85 341 119
rect 391 55 425 89
rect 570 73 604 107
rect 755 59 789 93
rect 859 68 893 102
rect 951 93 985 127
rect 1035 99 1069 133
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 119 427 153 461
rect 203 443 237 477
rect 203 375 237 409
rect 307 449 341 483
rect 307 381 341 415
rect 391 451 425 485
rect 391 383 425 417
rect 570 451 604 485
rect 755 451 789 485
rect 859 437 893 471
rect 859 334 893 368
rect 951 450 985 484
rect 951 330 985 364
rect 1035 441 1069 475
rect 1035 350 1069 384
<< poly >>
rect 609 366 673 376
rect 511 321 565 337
rect 609 332 623 366
rect 657 332 673 366
rect 609 322 673 332
rect 715 357 807 373
rect 715 323 763 357
rect 797 323 807 357
rect 511 287 521 321
rect 555 287 565 321
rect 715 307 807 323
rect 21 264 76 280
rect 21 230 32 264
rect 66 230 76 264
rect 21 214 76 230
rect 118 264 193 274
rect 511 271 565 287
rect 118 230 134 264
rect 168 230 193 264
rect 796 249 933 265
rect 118 220 193 230
rect 293 225 347 241
rect 293 191 303 225
rect 337 191 347 225
rect 293 175 347 191
rect 416 231 470 247
rect 416 197 426 231
rect 460 197 470 231
rect 796 215 806 249
rect 840 215 933 249
rect 416 183 470 197
rect 512 199 578 209
rect 796 199 933 215
rect 975 249 1034 265
rect 975 215 985 249
rect 1019 215 1034 249
rect 975 199 1034 215
rect 512 165 532 199
rect 566 165 578 199
rect 512 153 578 165
<< polycont >>
rect 623 332 657 366
rect 763 323 797 357
rect 521 287 555 321
rect 32 230 66 264
rect 134 230 168 264
rect 303 191 337 225
rect 426 197 460 231
rect 806 215 840 249
rect 985 215 1019 249
rect 532 165 566 199
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 35 477 69 493
rect 35 409 69 443
rect 103 461 169 527
rect 103 427 119 461
rect 153 427 169 461
rect 203 477 248 493
rect 391 485 449 527
rect 755 485 819 527
rect 237 443 248 477
rect 203 409 248 443
rect 69 375 156 393
rect 35 359 156 375
rect 17 264 66 325
rect 17 230 32 264
rect 17 197 66 230
rect 122 323 156 359
rect 122 280 156 289
rect 237 391 248 409
rect 203 357 214 375
rect 203 337 248 357
rect 286 449 307 483
rect 341 449 357 483
rect 286 415 357 449
rect 286 381 307 415
rect 341 381 357 415
rect 122 264 168 280
rect 122 230 134 264
rect 122 214 168 230
rect 122 161 156 214
rect 35 127 156 161
rect 35 119 69 127
rect 203 119 237 337
rect 286 333 357 381
rect 425 451 449 485
rect 549 451 570 485
rect 604 451 721 485
rect 391 417 449 451
rect 659 421 721 451
rect 789 451 819 485
rect 755 435 819 451
rect 859 471 908 487
rect 893 437 908 471
rect 659 418 724 421
rect 425 383 449 417
rect 678 417 724 418
rect 678 413 726 417
rect 678 409 729 413
rect 681 407 729 409
rect 686 402 729 407
rect 391 367 449 383
rect 489 391 556 401
rect 523 357 556 391
rect 286 299 423 333
rect 287 225 353 265
rect 287 191 303 225
rect 337 191 353 225
rect 389 247 423 299
rect 489 321 556 357
rect 489 287 521 321
rect 555 287 556 321
rect 489 271 556 287
rect 590 366 657 382
rect 590 332 623 366
rect 590 323 657 332
rect 624 312 657 323
rect 624 289 653 312
rect 691 290 729 402
rect 859 373 908 437
rect 763 368 908 373
rect 763 357 859 368
rect 797 334 859 357
rect 893 334 908 368
rect 797 323 908 334
rect 763 307 908 323
rect 944 484 1001 527
rect 944 450 951 484
rect 985 450 1001 484
rect 944 364 1001 450
rect 944 330 951 364
rect 985 330 1001 364
rect 1035 475 1087 491
rect 1069 441 1087 475
rect 1035 384 1087 441
rect 1069 350 1087 384
rect 1035 334 1087 350
rect 944 314 1001 330
rect 389 231 464 247
rect 389 197 426 231
rect 460 197 464 231
rect 590 208 653 289
rect 389 157 464 197
rect 35 69 69 85
rect 103 59 119 93
rect 153 59 169 93
rect 203 69 237 85
rect 302 153 464 157
rect 512 199 653 208
rect 512 165 532 199
rect 566 165 653 199
rect 302 123 423 153
rect 512 147 653 165
rect 687 265 729 290
rect 874 265 908 307
rect 687 249 840 265
rect 687 215 806 249
rect 687 199 840 215
rect 874 249 1019 265
rect 874 215 985 249
rect 874 199 1019 215
rect 302 119 341 123
rect 302 85 307 119
rect 687 107 721 199
rect 874 144 908 199
rect 1053 149 1087 334
rect 302 69 341 85
rect 103 17 169 59
rect 375 55 391 89
rect 425 55 441 89
rect 553 73 570 107
rect 604 73 721 107
rect 755 93 809 109
rect 375 17 441 55
rect 789 59 809 93
rect 755 17 809 59
rect 859 102 908 144
rect 893 68 908 102
rect 859 52 908 68
rect 951 127 996 143
rect 985 93 996 127
rect 951 17 996 93
rect 1035 133 1087 149
rect 1069 99 1087 133
rect 1035 83 1087 99
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 122 289 156 323
rect 214 375 237 391
rect 237 375 248 391
rect 214 357 248 375
rect 489 357 523 391
rect 590 289 624 323
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
<< metal1 >>
rect 0 561 1104 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 0 496 1104 527
rect 202 391 260 397
rect 202 357 214 391
rect 248 388 260 391
rect 477 391 535 397
rect 477 388 489 391
rect 248 360 489 388
rect 248 357 260 360
rect 202 351 260 357
rect 477 357 489 360
rect 523 357 535 391
rect 477 351 535 357
rect 110 323 168 329
rect 110 289 122 323
rect 156 320 168 323
rect 578 323 636 329
rect 578 320 590 323
rect 156 292 590 320
rect 156 289 168 292
rect 110 283 168 289
rect 578 289 590 292
rect 624 289 636 323
rect 578 283 636 289
rect 0 17 1104 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
rect 0 -48 1104 -17
<< labels >>
flabel locali s 305 221 339 255 0 FreeSans 200 0 0 0 D
port 1 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 GATE_N
port 2 nsew clock input
flabel locali s 1046 357 1080 391 0 FreeSans 200 0 0 0 Q
port 7 nsew signal output
flabel locali s 30 289 64 323 0 FreeSans 200 0 0 0 GATE_N
port 2 nsew clock input
flabel locali s 1046 425 1080 459 0 FreeSans 200 0 0 0 Q
port 7 nsew signal output
flabel locali s 1046 85 1080 119 0 FreeSans 200 0 0 0 Q
port 7 nsew signal output
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel nwell s 47 544 47 544 0 FreeSans 200 0 0 0 VPB
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel pwell s 47 0 47 0 0 FreeSans 200 0 0 0 VNB
rlabel comment s 0 0 0 0 4 dlxtn_1
rlabel metal1 s 0 -48 1104 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1104 592 1 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1104 544
string GDS_END 2859964
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2849362
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 27.600 0.000 
<< end >>
