magic
tech sky130A
magscale 1 2
timestamp 1681267127
<< locali >>
rect 243 689 559 708
rect 243 655 255 689
rect 289 655 337 689
rect 371 655 431 689
rect 465 655 513 689
rect 547 655 559 689
rect 243 617 559 655
rect 243 583 255 617
rect 289 583 337 617
rect 371 583 431 617
rect 465 583 513 617
rect 547 583 559 617
rect 243 569 559 583
rect 243 125 559 139
rect 243 91 255 125
rect 289 91 337 125
rect 371 91 431 125
rect 465 91 513 125
rect 547 91 559 125
rect 243 53 559 91
rect 243 19 255 53
rect 289 19 337 53
rect 371 19 431 53
rect 465 19 513 53
rect 547 19 559 53
rect 243 0 559 19
<< viali >>
rect 255 655 289 689
rect 337 655 371 689
rect 431 655 465 689
rect 513 655 547 689
rect 255 583 289 617
rect 337 583 371 617
rect 431 583 465 617
rect 513 583 547 617
rect 255 91 289 125
rect 337 91 371 125
rect 431 91 465 125
rect 513 91 547 125
rect 255 19 289 53
rect 337 19 371 53
rect 431 19 465 53
rect 513 19 547 53
<< obsli1 >>
rect 120 545 186 611
rect 616 545 682 611
rect 120 523 160 545
rect 642 523 682 545
rect 41 479 160 523
rect 41 445 60 479
rect 94 445 160 479
rect 41 407 160 445
rect 41 373 60 407
rect 94 373 160 407
rect 41 335 160 373
rect 41 301 60 335
rect 94 301 160 335
rect 41 263 160 301
rect 41 229 60 263
rect 94 229 160 263
rect 41 185 160 229
rect 212 185 246 523
rect 298 185 332 523
rect 384 185 418 523
rect 470 185 504 523
rect 556 185 590 523
rect 642 479 761 523
rect 642 445 708 479
rect 742 445 761 479
rect 642 407 761 445
rect 642 373 708 407
rect 742 373 761 407
rect 642 335 761 373
rect 642 301 708 335
rect 742 301 761 335
rect 642 263 761 301
rect 642 229 708 263
rect 742 229 761 263
rect 642 185 761 229
rect 120 163 160 185
rect 642 163 682 185
rect 120 97 186 163
rect 616 97 682 163
<< obsli1c >>
rect 60 445 94 479
rect 60 373 94 407
rect 60 301 94 335
rect 60 229 94 263
rect 708 445 742 479
rect 708 373 742 407
rect 708 301 742 335
rect 708 229 742 263
<< metal1 >>
rect 243 689 559 708
rect 243 655 255 689
rect 289 655 337 689
rect 371 655 431 689
rect 465 655 513 689
rect 547 655 559 689
rect 243 617 559 655
rect 243 583 255 617
rect 289 583 337 617
rect 371 583 431 617
rect 465 583 513 617
rect 547 583 559 617
rect 243 571 559 583
rect 41 479 100 507
rect 41 445 60 479
rect 94 445 100 479
rect 41 407 100 445
rect 41 373 60 407
rect 94 373 100 407
rect 41 335 100 373
rect 41 301 60 335
rect 94 301 100 335
rect 41 263 100 301
rect 41 229 60 263
rect 94 229 100 263
rect 41 201 100 229
rect 702 479 761 507
rect 702 445 708 479
rect 742 445 761 479
rect 702 407 761 445
rect 702 373 708 407
rect 742 373 761 407
rect 702 335 761 373
rect 702 301 708 335
rect 742 301 761 335
rect 702 263 761 301
rect 702 229 708 263
rect 742 229 761 263
rect 702 201 761 229
rect 243 125 559 137
rect 243 91 255 125
rect 289 91 337 125
rect 371 91 431 125
rect 465 91 513 125
rect 547 91 559 125
rect 243 53 559 91
rect 243 19 255 53
rect 289 19 337 53
rect 371 19 431 53
rect 465 19 513 53
rect 547 19 559 53
rect 243 0 559 19
<< obsm1 >>
rect 203 201 255 507
rect 289 201 341 507
rect 375 201 427 507
rect 461 201 513 507
rect 547 201 599 507
<< metal2 >>
rect 14 379 788 507
rect 14 201 788 329
<< labels >>
rlabel metal2 s 14 379 788 507 6 DRAIN
port 1 nsew
rlabel viali s 513 655 547 689 6 GATE
port 2 nsew
rlabel viali s 513 583 547 617 6 GATE
port 2 nsew
rlabel viali s 513 91 547 125 6 GATE
port 2 nsew
rlabel viali s 513 19 547 53 6 GATE
port 2 nsew
rlabel viali s 431 655 465 689 6 GATE
port 2 nsew
rlabel viali s 431 583 465 617 6 GATE
port 2 nsew
rlabel viali s 431 91 465 125 6 GATE
port 2 nsew
rlabel viali s 431 19 465 53 6 GATE
port 2 nsew
rlabel viali s 337 655 371 689 6 GATE
port 2 nsew
rlabel viali s 337 583 371 617 6 GATE
port 2 nsew
rlabel viali s 337 91 371 125 6 GATE
port 2 nsew
rlabel viali s 337 19 371 53 6 GATE
port 2 nsew
rlabel viali s 255 655 289 689 6 GATE
port 2 nsew
rlabel viali s 255 583 289 617 6 GATE
port 2 nsew
rlabel viali s 255 91 289 125 6 GATE
port 2 nsew
rlabel viali s 255 19 289 53 6 GATE
port 2 nsew
rlabel locali s 243 569 559 708 6 GATE
port 2 nsew
rlabel locali s 243 0 559 139 6 GATE
port 2 nsew
rlabel metal1 s 243 571 559 708 6 GATE
port 2 nsew
rlabel metal1 s 243 0 559 137 6 GATE
port 2 nsew
rlabel metal2 s 14 201 788 329 6 SOURCE
port 3 nsew
rlabel metal1 s 41 201 100 507 6 SUBSTRATE
port 4 nsew
rlabel metal1 s 702 201 761 507 6 SUBSTRATE
port 4 nsew
<< properties >>
string FIXED_BBOX 14 0 788 708
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 5530004
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 5515144
string device primitive
<< end >>
