magic
tech sky130A
magscale 1 2
timestamp 1681267127
use sky130_fd_io__com_pdpredrvr_pbiasv2  sky130_fd_io__com_pdpredrvr_pbiasv2_0
timestamp 1681267127
transform -1 0 20068 0 1 -2980
box 11368 2948 20000 5606
use sky130_fd_io__gpiov2_octl_mux  sky130_fd_io__gpiov2_octl_mux_0
timestamp 1681267127
transform 1 0 -1627 0 -1 3513
box 1191 1040 1945 3147
use sky130_fd_io__gpiov2_pdpredrvr_strong_nr2  sky130_fd_io__gpiov2_pdpredrvr_strong_nr2_0
timestamp 1681267127
transform 1 0 3465 0 -1 -331
box 4776 -2105 7725 -314
use sky130_fd_io__gpiov2_pdpredrvr_strong_nr3  sky130_fd_io__gpiov2_pdpredrvr_strong_nr3_0
timestamp 1681267127
transform -1 0 12458 0 1 3202
box 1191 -1273 2956 457
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_0
timestamp 1681267127
transform -1 0 -1117 0 -1 418
box 107 226 240 873
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_1
timestamp 1681267127
transform -1 0 -1117 0 -1 2582
box 107 226 240 873
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_0
timestamp 1681267127
transform 1 0 -1299 0 -1 418
box 107 226 460 873
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_1
timestamp 1681267127
transform 1 0 -1299 0 -1 2582
box 107 226 460 873
use sky130_fd_io__tk_em1o_cdns_5595914180880  sky130_fd_io__tk_em1o_cdns_5595914180880_0
timestamp 1681267127
transform 0 1 9429 1 0 1506
box 0 0 1 1
use sky130_fd_io__tk_em1o_cdns_5595914180880  sky130_fd_io__tk_em1o_cdns_5595914180880_1
timestamp 1681267127
transform 0 1 9829 -1 0 1806
box 0 0 1 1
use sky130_fd_io__tk_em1o_cdns_5595914180880  sky130_fd_io__tk_em1o_cdns_5595914180880_2
timestamp 1681267127
transform 1 0 9509 0 1 1481
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_5595914180882  sky130_fd_io__tk_em1s_cdns_5595914180882_0
timestamp 1681267127
transform -1 0 9455 0 -1 1675
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_5595914180882  sky130_fd_io__tk_em1s_cdns_5595914180882_1
timestamp 1681267127
transform 0 -1 9627 1 0 2680
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_5595914180882  sky130_fd_io__tk_em1s_cdns_5595914180882_2
timestamp 1681267127
transform -1 0 9518 0 1 1779
box 0 0 1 1
use sky130_fd_pr__model__nfet_highvoltage__example_55959141808139  sky130_fd_pr__model__nfet_highvoltage__example_55959141808139_0
timestamp 1681267127
transform 1 0 8867 0 1 1623
box -15 0 311 1
use sky130_fd_pr__model__nfet_highvoltage__example_55959141808183  sky130_fd_pr__model__nfet_highvoltage__example_55959141808183_0
timestamp 1681267127
transform 1 0 9247 0 1 1623
box -15 0 121 1
use sky130_fd_pr__model__nfet_highvoltage__example_55959141808369  sky130_fd_pr__model__nfet_highvoltage__example_55959141808369_0
timestamp 1681267127
transform 1 0 -1093 0 -1 596
box -1 0 121 1
use sky130_fd_pr__model__nfet_highvoltage__example_55959141808643  sky130_fd_pr__model__nfet_highvoltage__example_55959141808643_0
timestamp 1681267127
transform 1 0 -1373 0 -1 540
box -1 0 101 1
use sky130_fd_pr__model__pfet_highvoltage__example_55959141808141  sky130_fd_pr__model__pfet_highvoltage__example_55959141808141_0
timestamp 1681267127
transform 1 0 8867 0 -1 1363
box -15 0 -14 1
use sky130_fd_pr__model__pfet_highvoltage__example_55959141808141  sky130_fd_pr__model__pfet_highvoltage__example_55959141808141_1
timestamp 1681267127
transform -1 0 9163 0 -1 1363
box -15 0 -14 1
use sky130_fd_pr__model__pfet_highvoltage__example_55959141808184  sky130_fd_pr__model__pfet_highvoltage__example_55959141808184_0
timestamp 1681267127
transform 1 0 9247 0 -1 1363
box -15 0 121 1
use sky130_fd_pr__model__pfet_highvoltage__example_55959141808371  sky130_fd_pr__model__pfet_highvoltage__example_55959141808371_0
timestamp 1681267127
transform 1 0 -1093 0 -1 994
box -1 0 121 1
use sky130_fd_pr__model__pfet_highvoltage__example_55959141808371  sky130_fd_pr__model__pfet_highvoltage__example_55959141808371_1
timestamp 1681267127
transform 1 0 -1093 0 1 1062
box -1 0 121 1
use sky130_fd_pr__model__pfet_highvoltage__example_55959141808642  sky130_fd_pr__model__pfet_highvoltage__example_55959141808642_0
timestamp 1681267127
transform 1 0 -1373 0 -1 1394
box -1 0 101 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_0
timestamp 1681267127
transform 0 -1 -1228 -1 0 539
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_1
timestamp 1681267127
transform 0 -1 -1104 -1 0 539
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_2
timestamp 1681267127
transform 0 -1 -1104 1 0 1184
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_3
timestamp 1681267127
transform 0 -1 9222 -1 0 836
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_4
timestamp 1681267127
transform 1 0 9049 0 -1 1441
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_5
timestamp 1681267127
transform 1 0 8876 0 -1 1441
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_6
timestamp 1681267127
transform 0 1 9188 1 0 1741
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_7
timestamp 1681267127
transform 0 1 8808 1 0 1741
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_8
timestamp 1681267127
transform 1 0 8781 0 -1 1209
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_9
timestamp 1681267127
transform 1 0 6225 0 1 52
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_10
timestamp 1681267127
transform 1 0 9363 0 -1 1523
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_11
timestamp 1681267127
transform 0 -1 8726 -1 0 836
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_0
timestamp 1681267127
transform 1 0 9508 0 1 1779
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_1
timestamp 1681267127
transform -1 0 9881 0 1 2637
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_2
timestamp 1681267127
transform -1 0 9881 0 1 1779
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_3
timestamp 1681267127
transform -1 0 8848 0 1 1401
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_4
timestamp 1681267127
transform 1 0 6256 0 1 40
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_5
timestamp 1681267127
transform 1 0 6256 0 1 1073
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_6
timestamp 1681267127
transform 1 0 8172 0 1 406
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_7
timestamp 1681267127
transform 1 0 8628 0 1 876
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_8
timestamp 1681267127
transform 1 0 8628 0 1 1623
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_9
timestamp 1681267127
transform 1 0 6629 0 1 3027
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_10
timestamp 1681267127
transform 1 0 6705 0 1 1656
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_0
timestamp 1681267127
transform 0 -1 -999 -1 0 762
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_1
timestamp 1681267127
transform 0 1 8894 1 0 1395
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_2
timestamp 1681267127
transform 0 1 9070 1 0 1395
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_3
timestamp 1681267127
transform 0 1 9247 1 0 1395
box 0 0 1 1
<< properties >>
string GDS_END 7534196
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 7485506
<< end >>
